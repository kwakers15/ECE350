module multiplier(data_result, msb_data_result, data_resultRDY, data_exception, data_operandA, data_operandB, clock);
input [31:0] data_operandA, data_operandB;
input clock;
output [31:0] data_result, msb_data_result;
output data_resultRDY, data_exception;

assign data_resultRDY = 1'b1;

wire A0, A1, A2, A3, A4, A5, A6, A7, A8, A9, A10, A11, A12, A13, A14, A15, A16, A17, A18, A19, A20, A21, A22, A23, A24, A25, A26, A27, A28, A29, A30, A31;

assign A0 = data_operandA[0];
assign A1 = data_operandA[1];
assign A2 = data_operandA[2];
assign A3 = data_operandA[3];
assign A4 = data_operandA[4];
assign A5 = data_operandA[5];
assign A6 = data_operandA[6];
assign A7 = data_operandA[7];
assign A8 = data_operandA[8];
assign A9 = data_operandA[9];
assign A10 = data_operandA[10];
assign A11 = data_operandA[11];
assign A12 = data_operandA[12];
assign A13 = data_operandA[13];
assign A14 = data_operandA[14];
assign A15 = data_operandA[15];
assign A16 = data_operandA[16];
assign A17 = data_operandA[17];
assign A18 = data_operandA[18];
assign A19 = data_operandA[19];
assign A20 = data_operandA[20];
assign A21 = data_operandA[21];
assign A22 = data_operandA[22];
assign A23 = data_operandA[23];
assign A24 = data_operandA[24];
assign A25 = data_operandA[25];
assign A26 = data_operandA[26];
assign A27 = data_operandA[27];
assign A28 = data_operandA[28];
assign A29 = data_operandA[29];
assign A30 = data_operandA[30];
assign A31 = data_operandA[31];

wire B0, B1, B2, B3, B4, B5, B6, B7, B8, B9, B10, B11, B12, B13, B14, B15, B16, B17, B18, B19, B20, B21, B22, B23, B24, B25, B26, B27, B28, B29, B30, B31;

assign B0 = data_operandB[0];
assign B1 = data_operandB[1];
assign B2 = data_operandB[2];
assign B3 = data_operandB[3];
assign B4 = data_operandB[4];
assign B5 = data_operandB[5];
assign B6 = data_operandB[6];
assign B7 = data_operandB[7];
assign B8 = data_operandB[8];
assign B9 = data_operandB[9];
assign B10 = data_operandB[10];
assign B11 = data_operandB[11];
assign B12 = data_operandB[12];
assign B13 = data_operandB[13];
assign B14 = data_operandB[14];
assign B15 = data_operandB[15];
assign B16 = data_operandB[16];
assign B17 = data_operandB[17];
assign B18 = data_operandB[18];
assign B19 = data_operandB[19];
assign B20 = data_operandB[20];
assign B21 = data_operandB[21];
assign B22 = data_operandB[22];
assign B23 = data_operandB[23];
assign B24 = data_operandB[24];
assign B25 = data_operandB[25];
assign B26 = data_operandB[26];
assign B27 = data_operandB[27];
assign B28 = data_operandB[28];
assign B29 = data_operandB[29];
assign B30 = data_operandB[30];
assign B31 = data_operandB[31];

wire A0B0;

and A0B0_and(A0B0, A0, B0);

// bit position 0--------------------------------------------------


wire A1B0, A0B1;

and A1B0_and(A1B0, A1, B0);
and A0B1_and(A0B1, A0, B1);

// bit position 1--------------------------------------------------


wire A2B0, A1B1, A0B2;

and A2B0_and(A2B0, A2, B0);
and A1B1_and(A1B1, A1, B1);
and A0B2_and(A0B2, A0, B2);

// bit position 2--------------------------------------------------


wire A3B0, A2B1, A1B2, A0B3;

and A3B0_and(A3B0, A3, B0);
and A2B1_and(A2B1, A2, B1);
and A1B2_and(A1B2, A1, B2);
and A0B3_and(A0B3, A0, B3);

// bit position 3--------------------------------------------------


wire A4B0, A3B1, A2B2, A1B3, A0B4;

and A4B0_and(A4B0, A4, B0);
and A3B1_and(A3B1, A3, B1);
and A2B2_and(A2B2, A2, B2);
and A1B3_and(A1B3, A1, B3);
and A0B4_and(A0B4, A0, B4);

// bit position 4--------------------------------------------------


wire A5B0, A4B1, A3B2, A2B3, A1B4, A0B5;

and A5B0_and(A5B0, A5, B0);
and A4B1_and(A4B1, A4, B1);
and A3B2_and(A3B2, A3, B2);
and A2B3_and(A2B3, A2, B3);
and A1B4_and(A1B4, A1, B4);
and A0B5_and(A0B5, A0, B5);

// bit position 5--------------------------------------------------


wire A6B0, A5B1, A4B2, A3B3, A2B4, A1B5, A0B6;

and A6B0_and(A6B0, A6, B0);
and A5B1_and(A5B1, A5, B1);
and A4B2_and(A4B2, A4, B2);
and A3B3_and(A3B3, A3, B3);
and A2B4_and(A2B4, A2, B4);
and A1B5_and(A1B5, A1, B5);
and A0B6_and(A0B6, A0, B6);

// bit position 6--------------------------------------------------


wire A7B0, A6B1, A5B2, A4B3, A3B4, A2B5, A1B6, A0B7;

and A7B0_and(A7B0, A7, B0);
and A6B1_and(A6B1, A6, B1);
and A5B2_and(A5B2, A5, B2);
and A4B3_and(A4B3, A4, B3);
and A3B4_and(A3B4, A3, B4);
and A2B5_and(A2B5, A2, B5);
and A1B6_and(A1B6, A1, B6);
and A0B7_and(A0B7, A0, B7);

// bit position 7--------------------------------------------------


wire A8B0, A7B1, A6B2, A5B3, A4B4, A3B5, A2B6, A1B7, A0B8;

and A8B0_and(A8B0, A8, B0);
and A7B1_and(A7B1, A7, B1);
and A6B2_and(A6B2, A6, B2);
and A5B3_and(A5B3, A5, B3);
and A4B4_and(A4B4, A4, B4);
and A3B5_and(A3B5, A3, B5);
and A2B6_and(A2B6, A2, B6);
and A1B7_and(A1B7, A1, B7);
and A0B8_and(A0B8, A0, B8);

// bit position 8--------------------------------------------------


wire A9B0, A8B1, A7B2, A6B3, A5B4, A4B5, A3B6, A2B7, A1B8, A0B9;

and A9B0_and(A9B0, A9, B0);
and A8B1_and(A8B1, A8, B1);
and A7B2_and(A7B2, A7, B2);
and A6B3_and(A6B3, A6, B3);
and A5B4_and(A5B4, A5, B4);
and A4B5_and(A4B5, A4, B5);
and A3B6_and(A3B6, A3, B6);
and A2B7_and(A2B7, A2, B7);
and A1B8_and(A1B8, A1, B8);
and A0B9_and(A0B9, A0, B9);

// bit position 9--------------------------------------------------


wire A10B0, A9B1, A8B2, A7B3, A6B4, A5B5, A4B6, A3B7, A2B8, A1B9, A0B10;

and A10B0_and(A10B0, A10, B0);
and A9B1_and(A9B1, A9, B1);
and A8B2_and(A8B2, A8, B2);
and A7B3_and(A7B3, A7, B3);
and A6B4_and(A6B4, A6, B4);
and A5B5_and(A5B5, A5, B5);
and A4B6_and(A4B6, A4, B6);
and A3B7_and(A3B7, A3, B7);
and A2B8_and(A2B8, A2, B8);
and A1B9_and(A1B9, A1, B9);
and A0B10_and(A0B10, A0, B10);

// bit position 10--------------------------------------------------


wire A11B0, A10B1, A9B2, A8B3, A7B4, A6B5, A5B6, A4B7, A3B8, A2B9, A1B10, A0B11;

and A11B0_and(A11B0, A11, B0);
and A10B1_and(A10B1, A10, B1);
and A9B2_and(A9B2, A9, B2);
and A8B3_and(A8B3, A8, B3);
and A7B4_and(A7B4, A7, B4);
and A6B5_and(A6B5, A6, B5);
and A5B6_and(A5B6, A5, B6);
and A4B7_and(A4B7, A4, B7);
and A3B8_and(A3B8, A3, B8);
and A2B9_and(A2B9, A2, B9);
and A1B10_and(A1B10, A1, B10);
and A0B11_and(A0B11, A0, B11);

// bit position 11--------------------------------------------------


wire A12B0, A11B1, A10B2, A9B3, A8B4, A7B5, A6B6, A5B7, A4B8, A3B9, A2B10, A1B11, A0B12;

and A12B0_and(A12B0, A12, B0);
and A11B1_and(A11B1, A11, B1);
and A10B2_and(A10B2, A10, B2);
and A9B3_and(A9B3, A9, B3);
and A8B4_and(A8B4, A8, B4);
and A7B5_and(A7B5, A7, B5);
and A6B6_and(A6B6, A6, B6);
and A5B7_and(A5B7, A5, B7);
and A4B8_and(A4B8, A4, B8);
and A3B9_and(A3B9, A3, B9);
and A2B10_and(A2B10, A2, B10);
and A1B11_and(A1B11, A1, B11);
and A0B12_and(A0B12, A0, B12);

// bit position 12--------------------------------------------------


wire A13B0, A12B1, A11B2, A10B3, A9B4, A8B5, A7B6, A6B7, A5B8, A4B9, A3B10, A2B11, A1B12, A0B13;

and A13B0_and(A13B0, A13, B0);
and A12B1_and(A12B1, A12, B1);
and A11B2_and(A11B2, A11, B2);
and A10B3_and(A10B3, A10, B3);
and A9B4_and(A9B4, A9, B4);
and A8B5_and(A8B5, A8, B5);
and A7B6_and(A7B6, A7, B6);
and A6B7_and(A6B7, A6, B7);
and A5B8_and(A5B8, A5, B8);
and A4B9_and(A4B9, A4, B9);
and A3B10_and(A3B10, A3, B10);
and A2B11_and(A2B11, A2, B11);
and A1B12_and(A1B12, A1, B12);
and A0B13_and(A0B13, A0, B13);

// bit position 13--------------------------------------------------


wire A14B0, A13B1, A12B2, A11B3, A10B4, A9B5, A8B6, A7B7, A6B8, A5B9, A4B10, A3B11, A2B12, A1B13, A0B14;

and A14B0_and(A14B0, A14, B0);
and A13B1_and(A13B1, A13, B1);
and A12B2_and(A12B2, A12, B2);
and A11B3_and(A11B3, A11, B3);
and A10B4_and(A10B4, A10, B4);
and A9B5_and(A9B5, A9, B5);
and A8B6_and(A8B6, A8, B6);
and A7B7_and(A7B7, A7, B7);
and A6B8_and(A6B8, A6, B8);
and A5B9_and(A5B9, A5, B9);
and A4B10_and(A4B10, A4, B10);
and A3B11_and(A3B11, A3, B11);
and A2B12_and(A2B12, A2, B12);
and A1B13_and(A1B13, A1, B13);
and A0B14_and(A0B14, A0, B14);

// bit position 14--------------------------------------------------


wire A15B0, A14B1, A13B2, A12B3, A11B4, A10B5, A9B6, A8B7, A7B8, A6B9, A5B10, A4B11, A3B12, A2B13, A1B14, A0B15;

and A15B0_and(A15B0, A15, B0);
and A14B1_and(A14B1, A14, B1);
and A13B2_and(A13B2, A13, B2);
and A12B3_and(A12B3, A12, B3);
and A11B4_and(A11B4, A11, B4);
and A10B5_and(A10B5, A10, B5);
and A9B6_and(A9B6, A9, B6);
and A8B7_and(A8B7, A8, B7);
and A7B8_and(A7B8, A7, B8);
and A6B9_and(A6B9, A6, B9);
and A5B10_and(A5B10, A5, B10);
and A4B11_and(A4B11, A4, B11);
and A3B12_and(A3B12, A3, B12);
and A2B13_and(A2B13, A2, B13);
and A1B14_and(A1B14, A1, B14);
and A0B15_and(A0B15, A0, B15);

// bit position 15--------------------------------------------------


wire A16B0, A15B1, A14B2, A13B3, A12B4, A11B5, A10B6, A9B7, A8B8, A7B9, A6B10, A5B11, A4B12, A3B13, A2B14, A1B15, A0B16;

and A16B0_and(A16B0, A16, B0);
and A15B1_and(A15B1, A15, B1);
and A14B2_and(A14B2, A14, B2);
and A13B3_and(A13B3, A13, B3);
and A12B4_and(A12B4, A12, B4);
and A11B5_and(A11B5, A11, B5);
and A10B6_and(A10B6, A10, B6);
and A9B7_and(A9B7, A9, B7);
and A8B8_and(A8B8, A8, B8);
and A7B9_and(A7B9, A7, B9);
and A6B10_and(A6B10, A6, B10);
and A5B11_and(A5B11, A5, B11);
and A4B12_and(A4B12, A4, B12);
and A3B13_and(A3B13, A3, B13);
and A2B14_and(A2B14, A2, B14);
and A1B15_and(A1B15, A1, B15);
and A0B16_and(A0B16, A0, B16);

// bit position 16--------------------------------------------------


wire A17B0, A16B1, A15B2, A14B3, A13B4, A12B5, A11B6, A10B7, A9B8, A8B9, A7B10, A6B11, A5B12, A4B13, A3B14, A2B15, A1B16, A0B17;

and A17B0_and(A17B0, A17, B0);
and A16B1_and(A16B1, A16, B1);
and A15B2_and(A15B2, A15, B2);
and A14B3_and(A14B3, A14, B3);
and A13B4_and(A13B4, A13, B4);
and A12B5_and(A12B5, A12, B5);
and A11B6_and(A11B6, A11, B6);
and A10B7_and(A10B7, A10, B7);
and A9B8_and(A9B8, A9, B8);
and A8B9_and(A8B9, A8, B9);
and A7B10_and(A7B10, A7, B10);
and A6B11_and(A6B11, A6, B11);
and A5B12_and(A5B12, A5, B12);
and A4B13_and(A4B13, A4, B13);
and A3B14_and(A3B14, A3, B14);
and A2B15_and(A2B15, A2, B15);
and A1B16_and(A1B16, A1, B16);
and A0B17_and(A0B17, A0, B17);

// bit position 17--------------------------------------------------


wire A18B0, A17B1, A16B2, A15B3, A14B4, A13B5, A12B6, A11B7, A10B8, A9B9, A8B10, A7B11, A6B12, A5B13, A4B14, A3B15, A2B16, A1B17, A0B18;

and A18B0_and(A18B0, A18, B0);
and A17B1_and(A17B1, A17, B1);
and A16B2_and(A16B2, A16, B2);
and A15B3_and(A15B3, A15, B3);
and A14B4_and(A14B4, A14, B4);
and A13B5_and(A13B5, A13, B5);
and A12B6_and(A12B6, A12, B6);
and A11B7_and(A11B7, A11, B7);
and A10B8_and(A10B8, A10, B8);
and A9B9_and(A9B9, A9, B9);
and A8B10_and(A8B10, A8, B10);
and A7B11_and(A7B11, A7, B11);
and A6B12_and(A6B12, A6, B12);
and A5B13_and(A5B13, A5, B13);
and A4B14_and(A4B14, A4, B14);
and A3B15_and(A3B15, A3, B15);
and A2B16_and(A2B16, A2, B16);
and A1B17_and(A1B17, A1, B17);
and A0B18_and(A0B18, A0, B18);

// bit position 18--------------------------------------------------


wire A19B0, A18B1, A17B2, A16B3, A15B4, A14B5, A13B6, A12B7, A11B8, A10B9, A9B10, A8B11, A7B12, A6B13, A5B14, A4B15, A3B16, A2B17, A1B18, A0B19;

and A19B0_and(A19B0, A19, B0);
and A18B1_and(A18B1, A18, B1);
and A17B2_and(A17B2, A17, B2);
and A16B3_and(A16B3, A16, B3);
and A15B4_and(A15B4, A15, B4);
and A14B5_and(A14B5, A14, B5);
and A13B6_and(A13B6, A13, B6);
and A12B7_and(A12B7, A12, B7);
and A11B8_and(A11B8, A11, B8);
and A10B9_and(A10B9, A10, B9);
and A9B10_and(A9B10, A9, B10);
and A8B11_and(A8B11, A8, B11);
and A7B12_and(A7B12, A7, B12);
and A6B13_and(A6B13, A6, B13);
and A5B14_and(A5B14, A5, B14);
and A4B15_and(A4B15, A4, B15);
and A3B16_and(A3B16, A3, B16);
and A2B17_and(A2B17, A2, B17);
and A1B18_and(A1B18, A1, B18);
and A0B19_and(A0B19, A0, B19);

// bit position 19--------------------------------------------------


wire A20B0, A19B1, A18B2, A17B3, A16B4, A15B5, A14B6, A13B7, A12B8, A11B9, A10B10, A9B11, A8B12, A7B13, A6B14, A5B15, A4B16, A3B17, A2B18, A1B19, A0B20;

and A20B0_and(A20B0, A20, B0);
and A19B1_and(A19B1, A19, B1);
and A18B2_and(A18B2, A18, B2);
and A17B3_and(A17B3, A17, B3);
and A16B4_and(A16B4, A16, B4);
and A15B5_and(A15B5, A15, B5);
and A14B6_and(A14B6, A14, B6);
and A13B7_and(A13B7, A13, B7);
and A12B8_and(A12B8, A12, B8);
and A11B9_and(A11B9, A11, B9);
and A10B10_and(A10B10, A10, B10);
and A9B11_and(A9B11, A9, B11);
and A8B12_and(A8B12, A8, B12);
and A7B13_and(A7B13, A7, B13);
and A6B14_and(A6B14, A6, B14);
and A5B15_and(A5B15, A5, B15);
and A4B16_and(A4B16, A4, B16);
and A3B17_and(A3B17, A3, B17);
and A2B18_and(A2B18, A2, B18);
and A1B19_and(A1B19, A1, B19);
and A0B20_and(A0B20, A0, B20);

// bit position 20--------------------------------------------------


wire A21B0, A20B1, A19B2, A18B3, A17B4, A16B5, A15B6, A14B7, A13B8, A12B9, A11B10, A10B11, A9B12, A8B13, A7B14, A6B15, A5B16, A4B17, A3B18, A2B19, A1B20, A0B21;

and A21B0_and(A21B0, A21, B0);
and A20B1_and(A20B1, A20, B1);
and A19B2_and(A19B2, A19, B2);
and A18B3_and(A18B3, A18, B3);
and A17B4_and(A17B4, A17, B4);
and A16B5_and(A16B5, A16, B5);
and A15B6_and(A15B6, A15, B6);
and A14B7_and(A14B7, A14, B7);
and A13B8_and(A13B8, A13, B8);
and A12B9_and(A12B9, A12, B9);
and A11B10_and(A11B10, A11, B10);
and A10B11_and(A10B11, A10, B11);
and A9B12_and(A9B12, A9, B12);
and A8B13_and(A8B13, A8, B13);
and A7B14_and(A7B14, A7, B14);
and A6B15_and(A6B15, A6, B15);
and A5B16_and(A5B16, A5, B16);
and A4B17_and(A4B17, A4, B17);
and A3B18_and(A3B18, A3, B18);
and A2B19_and(A2B19, A2, B19);
and A1B20_and(A1B20, A1, B20);
and A0B21_and(A0B21, A0, B21);

// bit position 21--------------------------------------------------


wire A22B0, A21B1, A20B2, A19B3, A18B4, A17B5, A16B6, A15B7, A14B8, A13B9, A12B10, A11B11, A10B12, A9B13, A8B14, A7B15, A6B16, A5B17, A4B18, A3B19, A2B20, A1B21, A0B22;

and A22B0_and(A22B0, A22, B0);
and A21B1_and(A21B1, A21, B1);
and A20B2_and(A20B2, A20, B2);
and A19B3_and(A19B3, A19, B3);
and A18B4_and(A18B4, A18, B4);
and A17B5_and(A17B5, A17, B5);
and A16B6_and(A16B6, A16, B6);
and A15B7_and(A15B7, A15, B7);
and A14B8_and(A14B8, A14, B8);
and A13B9_and(A13B9, A13, B9);
and A12B10_and(A12B10, A12, B10);
and A11B11_and(A11B11, A11, B11);
and A10B12_and(A10B12, A10, B12);
and A9B13_and(A9B13, A9, B13);
and A8B14_and(A8B14, A8, B14);
and A7B15_and(A7B15, A7, B15);
and A6B16_and(A6B16, A6, B16);
and A5B17_and(A5B17, A5, B17);
and A4B18_and(A4B18, A4, B18);
and A3B19_and(A3B19, A3, B19);
and A2B20_and(A2B20, A2, B20);
and A1B21_and(A1B21, A1, B21);
and A0B22_and(A0B22, A0, B22);

// bit position 22--------------------------------------------------


wire A23B0, A22B1, A21B2, A20B3, A19B4, A18B5, A17B6, A16B7, A15B8, A14B9, A13B10, A12B11, A11B12, A10B13, A9B14, A8B15, A7B16, A6B17, A5B18, A4B19, A3B20, A2B21, A1B22, A0B23;

and A23B0_and(A23B0, A23, B0);
and A22B1_and(A22B1, A22, B1);
and A21B2_and(A21B2, A21, B2);
and A20B3_and(A20B3, A20, B3);
and A19B4_and(A19B4, A19, B4);
and A18B5_and(A18B5, A18, B5);
and A17B6_and(A17B6, A17, B6);
and A16B7_and(A16B7, A16, B7);
and A15B8_and(A15B8, A15, B8);
and A14B9_and(A14B9, A14, B9);
and A13B10_and(A13B10, A13, B10);
and A12B11_and(A12B11, A12, B11);
and A11B12_and(A11B12, A11, B12);
and A10B13_and(A10B13, A10, B13);
and A9B14_and(A9B14, A9, B14);
and A8B15_and(A8B15, A8, B15);
and A7B16_and(A7B16, A7, B16);
and A6B17_and(A6B17, A6, B17);
and A5B18_and(A5B18, A5, B18);
and A4B19_and(A4B19, A4, B19);
and A3B20_and(A3B20, A3, B20);
and A2B21_and(A2B21, A2, B21);
and A1B22_and(A1B22, A1, B22);
and A0B23_and(A0B23, A0, B23);

// bit position 23--------------------------------------------------


wire A24B0, A23B1, A22B2, A21B3, A20B4, A19B5, A18B6, A17B7, A16B8, A15B9, A14B10, A13B11, A12B12, A11B13, A10B14, A9B15, A8B16, A7B17, A6B18, A5B19, A4B20, A3B21, A2B22, A1B23, A0B24;

and A24B0_and(A24B0, A24, B0);
and A23B1_and(A23B1, A23, B1);
and A22B2_and(A22B2, A22, B2);
and A21B3_and(A21B3, A21, B3);
and A20B4_and(A20B4, A20, B4);
and A19B5_and(A19B5, A19, B5);
and A18B6_and(A18B6, A18, B6);
and A17B7_and(A17B7, A17, B7);
and A16B8_and(A16B8, A16, B8);
and A15B9_and(A15B9, A15, B9);
and A14B10_and(A14B10, A14, B10);
and A13B11_and(A13B11, A13, B11);
and A12B12_and(A12B12, A12, B12);
and A11B13_and(A11B13, A11, B13);
and A10B14_and(A10B14, A10, B14);
and A9B15_and(A9B15, A9, B15);
and A8B16_and(A8B16, A8, B16);
and A7B17_and(A7B17, A7, B17);
and A6B18_and(A6B18, A6, B18);
and A5B19_and(A5B19, A5, B19);
and A4B20_and(A4B20, A4, B20);
and A3B21_and(A3B21, A3, B21);
and A2B22_and(A2B22, A2, B22);
and A1B23_and(A1B23, A1, B23);
and A0B24_and(A0B24, A0, B24);

// bit position 24--------------------------------------------------


wire A25B0, A24B1, A23B2, A22B3, A21B4, A20B5, A19B6, A18B7, A17B8, A16B9, A15B10, A14B11, A13B12, A12B13, A11B14, A10B15, A9B16, A8B17, A7B18, A6B19, A5B20, A4B21, A3B22, A2B23, A1B24, A0B25;

and A25B0_and(A25B0, A25, B0);
and A24B1_and(A24B1, A24, B1);
and A23B2_and(A23B2, A23, B2);
and A22B3_and(A22B3, A22, B3);
and A21B4_and(A21B4, A21, B4);
and A20B5_and(A20B5, A20, B5);
and A19B6_and(A19B6, A19, B6);
and A18B7_and(A18B7, A18, B7);
and A17B8_and(A17B8, A17, B8);
and A16B9_and(A16B9, A16, B9);
and A15B10_and(A15B10, A15, B10);
and A14B11_and(A14B11, A14, B11);
and A13B12_and(A13B12, A13, B12);
and A12B13_and(A12B13, A12, B13);
and A11B14_and(A11B14, A11, B14);
and A10B15_and(A10B15, A10, B15);
and A9B16_and(A9B16, A9, B16);
and A8B17_and(A8B17, A8, B17);
and A7B18_and(A7B18, A7, B18);
and A6B19_and(A6B19, A6, B19);
and A5B20_and(A5B20, A5, B20);
and A4B21_and(A4B21, A4, B21);
and A3B22_and(A3B22, A3, B22);
and A2B23_and(A2B23, A2, B23);
and A1B24_and(A1B24, A1, B24);
and A0B25_and(A0B25, A0, B25);

// bit position 25--------------------------------------------------


wire A26B0, A25B1, A24B2, A23B3, A22B4, A21B5, A20B6, A19B7, A18B8, A17B9, A16B10, A15B11, A14B12, A13B13, A12B14, A11B15, A10B16, A9B17, A8B18, A7B19, A6B20, A5B21, A4B22, A3B23, A2B24, A1B25, A0B26;

and A26B0_and(A26B0, A26, B0);
and A25B1_and(A25B1, A25, B1);
and A24B2_and(A24B2, A24, B2);
and A23B3_and(A23B3, A23, B3);
and A22B4_and(A22B4, A22, B4);
and A21B5_and(A21B5, A21, B5);
and A20B6_and(A20B6, A20, B6);
and A19B7_and(A19B7, A19, B7);
and A18B8_and(A18B8, A18, B8);
and A17B9_and(A17B9, A17, B9);
and A16B10_and(A16B10, A16, B10);
and A15B11_and(A15B11, A15, B11);
and A14B12_and(A14B12, A14, B12);
and A13B13_and(A13B13, A13, B13);
and A12B14_and(A12B14, A12, B14);
and A11B15_and(A11B15, A11, B15);
and A10B16_and(A10B16, A10, B16);
and A9B17_and(A9B17, A9, B17);
and A8B18_and(A8B18, A8, B18);
and A7B19_and(A7B19, A7, B19);
and A6B20_and(A6B20, A6, B20);
and A5B21_and(A5B21, A5, B21);
and A4B22_and(A4B22, A4, B22);
and A3B23_and(A3B23, A3, B23);
and A2B24_and(A2B24, A2, B24);
and A1B25_and(A1B25, A1, B25);
and A0B26_and(A0B26, A0, B26);

// bit position 26--------------------------------------------------


wire A27B0, A26B1, A25B2, A24B3, A23B4, A22B5, A21B6, A20B7, A19B8, A18B9, A17B10, A16B11, A15B12, A14B13, A13B14, A12B15, A11B16, A10B17, A9B18, A8B19, A7B20, A6B21, A5B22, A4B23, A3B24, A2B25, A1B26, A0B27;

and A27B0_and(A27B0, A27, B0);
and A26B1_and(A26B1, A26, B1);
and A25B2_and(A25B2, A25, B2);
and A24B3_and(A24B3, A24, B3);
and A23B4_and(A23B4, A23, B4);
and A22B5_and(A22B5, A22, B5);
and A21B6_and(A21B6, A21, B6);
and A20B7_and(A20B7, A20, B7);
and A19B8_and(A19B8, A19, B8);
and A18B9_and(A18B9, A18, B9);
and A17B10_and(A17B10, A17, B10);
and A16B11_and(A16B11, A16, B11);
and A15B12_and(A15B12, A15, B12);
and A14B13_and(A14B13, A14, B13);
and A13B14_and(A13B14, A13, B14);
and A12B15_and(A12B15, A12, B15);
and A11B16_and(A11B16, A11, B16);
and A10B17_and(A10B17, A10, B17);
and A9B18_and(A9B18, A9, B18);
and A8B19_and(A8B19, A8, B19);
and A7B20_and(A7B20, A7, B20);
and A6B21_and(A6B21, A6, B21);
and A5B22_and(A5B22, A5, B22);
and A4B23_and(A4B23, A4, B23);
and A3B24_and(A3B24, A3, B24);
and A2B25_and(A2B25, A2, B25);
and A1B26_and(A1B26, A1, B26);
and A0B27_and(A0B27, A0, B27);

// bit position 27--------------------------------------------------


wire A28B0, A27B1, A26B2, A25B3, A24B4, A23B5, A22B6, A21B7, A20B8, A19B9, A18B10, A17B11, A16B12, A15B13, A14B14, A13B15, A12B16, A11B17, A10B18, A9B19, A8B20, A7B21, A6B22, A5B23, A4B24, A3B25, A2B26, A1B27, A0B28;

and A28B0_and(A28B0, A28, B0);
and A27B1_and(A27B1, A27, B1);
and A26B2_and(A26B2, A26, B2);
and A25B3_and(A25B3, A25, B3);
and A24B4_and(A24B4, A24, B4);
and A23B5_and(A23B5, A23, B5);
and A22B6_and(A22B6, A22, B6);
and A21B7_and(A21B7, A21, B7);
and A20B8_and(A20B8, A20, B8);
and A19B9_and(A19B9, A19, B9);
and A18B10_and(A18B10, A18, B10);
and A17B11_and(A17B11, A17, B11);
and A16B12_and(A16B12, A16, B12);
and A15B13_and(A15B13, A15, B13);
and A14B14_and(A14B14, A14, B14);
and A13B15_and(A13B15, A13, B15);
and A12B16_and(A12B16, A12, B16);
and A11B17_and(A11B17, A11, B17);
and A10B18_and(A10B18, A10, B18);
and A9B19_and(A9B19, A9, B19);
and A8B20_and(A8B20, A8, B20);
and A7B21_and(A7B21, A7, B21);
and A6B22_and(A6B22, A6, B22);
and A5B23_and(A5B23, A5, B23);
and A4B24_and(A4B24, A4, B24);
and A3B25_and(A3B25, A3, B25);
and A2B26_and(A2B26, A2, B26);
and A1B27_and(A1B27, A1, B27);
and A0B28_and(A0B28, A0, B28);

// bit position 28--------------------------------------------------


wire A29B0, A28B1, A27B2, A26B3, A25B4, A24B5, A23B6, A22B7, A21B8, A20B9, A19B10, A18B11, A17B12, A16B13, A15B14, A14B15, A13B16, A12B17, A11B18, A10B19, A9B20, A8B21, A7B22, A6B23, A5B24, A4B25, A3B26, A2B27, A1B28, A0B29;

and A29B0_and(A29B0, A29, B0);
and A28B1_and(A28B1, A28, B1);
and A27B2_and(A27B2, A27, B2);
and A26B3_and(A26B3, A26, B3);
and A25B4_and(A25B4, A25, B4);
and A24B5_and(A24B5, A24, B5);
and A23B6_and(A23B6, A23, B6);
and A22B7_and(A22B7, A22, B7);
and A21B8_and(A21B8, A21, B8);
and A20B9_and(A20B9, A20, B9);
and A19B10_and(A19B10, A19, B10);
and A18B11_and(A18B11, A18, B11);
and A17B12_and(A17B12, A17, B12);
and A16B13_and(A16B13, A16, B13);
and A15B14_and(A15B14, A15, B14);
and A14B15_and(A14B15, A14, B15);
and A13B16_and(A13B16, A13, B16);
and A12B17_and(A12B17, A12, B17);
and A11B18_and(A11B18, A11, B18);
and A10B19_and(A10B19, A10, B19);
and A9B20_and(A9B20, A9, B20);
and A8B21_and(A8B21, A8, B21);
and A7B22_and(A7B22, A7, B22);
and A6B23_and(A6B23, A6, B23);
and A5B24_and(A5B24, A5, B24);
and A4B25_and(A4B25, A4, B25);
and A3B26_and(A3B26, A3, B26);
and A2B27_and(A2B27, A2, B27);
and A1B28_and(A1B28, A1, B28);
and A0B29_and(A0B29, A0, B29);

// bit position 29--------------------------------------------------


wire A30B0, A29B1, A28B2, A27B3, A26B4, A25B5, A24B6, A23B7, A22B8, A21B9, A20B10, A19B11, A18B12, A17B13, A16B14, A15B15, A14B16, A13B17, A12B18, A11B19, A10B20, A9B21, A8B22, A7B23, A6B24, A5B25, A4B26, A3B27, A2B28, A1B29, A0B30;

and A30B0_and(A30B0, A30, B0);
and A29B1_and(A29B1, A29, B1);
and A28B2_and(A28B2, A28, B2);
and A27B3_and(A27B3, A27, B3);
and A26B4_and(A26B4, A26, B4);
and A25B5_and(A25B5, A25, B5);
and A24B6_and(A24B6, A24, B6);
and A23B7_and(A23B7, A23, B7);
and A22B8_and(A22B8, A22, B8);
and A21B9_and(A21B9, A21, B9);
and A20B10_and(A20B10, A20, B10);
and A19B11_and(A19B11, A19, B11);
and A18B12_and(A18B12, A18, B12);
and A17B13_and(A17B13, A17, B13);
and A16B14_and(A16B14, A16, B14);
and A15B15_and(A15B15, A15, B15);
and A14B16_and(A14B16, A14, B16);
and A13B17_and(A13B17, A13, B17);
and A12B18_and(A12B18, A12, B18);
and A11B19_and(A11B19, A11, B19);
and A10B20_and(A10B20, A10, B20);
and A9B21_and(A9B21, A9, B21);
and A8B22_and(A8B22, A8, B22);
and A7B23_and(A7B23, A7, B23);
and A6B24_and(A6B24, A6, B24);
and A5B25_and(A5B25, A5, B25);
and A4B26_and(A4B26, A4, B26);
and A3B27_and(A3B27, A3, B27);
and A2B28_and(A2B28, A2, B28);
and A1B29_and(A1B29, A1, B29);
and A0B30_and(A0B30, A0, B30);

// bit position 30--------------------------------------------------


wire A31B0, A30B1, A29B2, A28B3, A27B4, A26B5, A25B6, A24B7, A23B8, A22B9, A21B10, A20B11, A19B12, A18B13, A17B14, A16B15, A15B16, A14B17, A13B18, A12B19, A11B20, A10B21, A9B22, A8B23, A7B24, A6B25, A5B26, A4B27, A3B28, A2B29, A1B30, A0B31;

and A31B0_and(A31B0, A31, B0);
and A30B1_and(A30B1, A30, B1);
and A29B2_and(A29B2, A29, B2);
and A28B3_and(A28B3, A28, B3);
and A27B4_and(A27B4, A27, B4);
and A26B5_and(A26B5, A26, B5);
and A25B6_and(A25B6, A25, B6);
and A24B7_and(A24B7, A24, B7);
and A23B8_and(A23B8, A23, B8);
and A22B9_and(A22B9, A22, B9);
and A21B10_and(A21B10, A21, B10);
and A20B11_and(A20B11, A20, B11);
and A19B12_and(A19B12, A19, B12);
and A18B13_and(A18B13, A18, B13);
and A17B14_and(A17B14, A17, B14);
and A16B15_and(A16B15, A16, B15);
and A15B16_and(A15B16, A15, B16);
and A14B17_and(A14B17, A14, B17);
and A13B18_and(A13B18, A13, B18);
and A12B19_and(A12B19, A12, B19);
and A11B20_and(A11B20, A11, B20);
and A10B21_and(A10B21, A10, B21);
and A9B22_and(A9B22, A9, B22);
and A8B23_and(A8B23, A8, B23);
and A7B24_and(A7B24, A7, B24);
and A6B25_and(A6B25, A6, B25);
and A5B26_and(A5B26, A5, B26);
and A4B27_and(A4B27, A4, B27);
and A3B28_and(A3B28, A3, B28);
and A2B29_and(A2B29, A2, B29);
and A1B30_and(A1B30, A1, B30);
and A0B31_and(A0B31, A0, B31);

// bit position 31--------------------------------------------------

wire A31B1, A30B2, A29B3, A28B4, A27B5, A26B6, A25B7, A24B8, A23B9, A22B10, A21B11, A20B12, A19B13, A18B14, A17B15, A16B16, A15B17, A14B18, A13B19, A12B20, A11B21, A10B22, A9B23, A8B24, A7B25, A6B26, A5B27, A4B28, A3B29, A2B30, A1B31;

and A31B1_and(A31B1, A31, B1);
and A30B2_and(A30B2, A30, B2);
and A29B3_and(A29B3, A29, B3);
and A28B4_and(A28B4, A28, B4);
and A27B5_and(A27B5, A27, B5);
and A26B6_and(A26B6, A26, B6);
and A25B7_and(A25B7, A25, B7);
and A24B8_and(A24B8, A24, B8);
and A23B9_and(A23B9, A23, B9);
and A22B10_and(A22B10, A22, B10);
and A21B11_and(A21B11, A21, B11);
and A20B12_and(A20B12, A20, B12);
and A19B13_and(A19B13, A19, B13);
and A18B14_and(A18B14, A18, B14);
and A17B15_and(A17B15, A17, B15);
and A16B16_and(A16B16, A16, B16);
and A15B17_and(A15B17, A15, B17);
and A14B18_and(A14B18, A14, B18);
and A13B19_and(A13B19, A13, B19);
and A12B20_and(A12B20, A12, B20);
and A11B21_and(A11B21, A11, B21);
and A10B22_and(A10B22, A10, B22);
and A9B23_and(A9B23, A9, B23);
and A8B24_and(A8B24, A8, B24);
and A7B25_and(A7B25, A7, B25);
and A6B26_and(A6B26, A6, B26);
and A5B27_and(A5B27, A5, B27);
and A4B28_and(A4B28, A4, B28);
and A3B29_and(A3B29, A3, B29);
and A2B30_and(A2B30, A2, B30);
and A1B31_and(A1B31, A1, B31);

// bit position 32------------------------------------------------------------

wire A31B2, A30B3, A29B4, A28B5, A27B6, A26B7, A25B8, A24B9, A23B10, A22B11, A21B12, A20B13, A19B14, A18B15, A17B16, A16B17, A15B18, A14B19, A13B20, A12B21, A11B22, A10B23, A9B24, A8B25, A7B26, A6B27, A5B28, A4B29, A3B30, A2B31;

and A31B2_and(A31B2, A31, B2);
and A30B3_and(A30B3, A30, B3);
and A29B4_and(A29B4, A29, B4);
and A28B5_and(A28B5, A28, B5);
and A27B6_and(A27B6, A27, B6);
and A26B7_and(A26B7, A26, B7);
and A25B8_and(A25B8, A25, B8);
and A24B9_and(A24B9, A24, B9);
and A23B10_and(A23B10, A23, B10);
and A22B11_and(A22B11, A22, B11);
and A21B12_and(A21B12, A21, B12);
and A20B13_and(A20B13, A20, B13);
and A19B14_and(A19B14, A19, B14);
and A18B15_and(A18B15, A18, B15);
and A17B16_and(A17B16, A17, B16);
and A16B17_and(A16B17, A16, B17);
and A15B18_and(A15B18, A15, B18);
and A14B19_and(A14B19, A14, B19);
and A13B20_and(A13B20, A13, B20);
and A12B21_and(A12B21, A12, B21);
and A11B22_and(A11B22, A11, B22);
and A10B23_and(A10B23, A10, B23);
and A9B24_and(A9B24, A9, B24);
and A8B25_and(A8B25, A8, B25);
and A7B26_and(A7B26, A7, B26);
and A6B27_and(A6B27, A6, B27);
and A5B28_and(A5B28, A5, B28);
and A4B29_and(A4B29, A4, B29);
and A3B30_and(A3B30, A3, B30);
and A2B31_and(A2B31, A2, B31);

// bit position 33------------------------------------------------------------

wire A31B3, A30B4, A29B5, A28B6, A27B7, A26B8, A25B9, A24B10, A23B11, A22B12, A21B13, A20B14, A19B15, A18B16, A17B17, A16B18, A15B19, A14B20, A13B21, A12B22, A11B23, A10B24, A9B25, A8B26, A7B27, A6B28, A5B29, A4B30, A3B31;

and A31B3_and(A31B3, A31, B3);
and A30B4_and(A30B4, A30, B4);
and A29B5_and(A29B5, A29, B5);
and A28B6_and(A28B6, A28, B6);
and A27B7_and(A27B7, A27, B7);
and A26B8_and(A26B8, A26, B8);
and A25B9_and(A25B9, A25, B9);
and A24B10_and(A24B10, A24, B10);
and A23B11_and(A23B11, A23, B11);
and A22B12_and(A22B12, A22, B12);
and A21B13_and(A21B13, A21, B13);
and A20B14_and(A20B14, A20, B14);
and A19B15_and(A19B15, A19, B15);
and A18B16_and(A18B16, A18, B16);
and A17B17_and(A17B17, A17, B17);
and A16B18_and(A16B18, A16, B18);
and A15B19_and(A15B19, A15, B19);
and A14B20_and(A14B20, A14, B20);
and A13B21_and(A13B21, A13, B21);
and A12B22_and(A12B22, A12, B22);
and A11B23_and(A11B23, A11, B23);
and A10B24_and(A10B24, A10, B24);
and A9B25_and(A9B25, A9, B25);
and A8B26_and(A8B26, A8, B26);
and A7B27_and(A7B27, A7, B27);
and A6B28_and(A6B28, A6, B28);
and A5B29_and(A5B29, A5, B29);
and A4B30_and(A4B30, A4, B30);
and A3B31_and(A3B31, A3, B31);

// bit position 34------------------------------------------------------------

wire A31B4, A30B5, A29B6, A28B7, A27B8, A26B9, A25B10, A24B11, A23B12, A22B13, A21B14, A20B15, A19B16, A18B17, A17B18, A16B19, A15B20, A14B21, A13B22, A12B23, A11B24, A10B25, A9B26, A8B27, A7B28, A6B29, A5B30, A4B31;

and A31B4_and(A31B4, A31, B4);
and A30B5_and(A30B5, A30, B5);
and A29B6_and(A29B6, A29, B6);
and A28B7_and(A28B7, A28, B7);
and A27B8_and(A27B8, A27, B8);
and A26B9_and(A26B9, A26, B9);
and A25B10_and(A25B10, A25, B10);
and A24B11_and(A24B11, A24, B11);
and A23B12_and(A23B12, A23, B12);
and A22B13_and(A22B13, A22, B13);
and A21B14_and(A21B14, A21, B14);
and A20B15_and(A20B15, A20, B15);
and A19B16_and(A19B16, A19, B16);
and A18B17_and(A18B17, A18, B17);
and A17B18_and(A17B18, A17, B18);
and A16B19_and(A16B19, A16, B19);
and A15B20_and(A15B20, A15, B20);
and A14B21_and(A14B21, A14, B21);
and A13B22_and(A13B22, A13, B22);
and A12B23_and(A12B23, A12, B23);
and A11B24_and(A11B24, A11, B24);
and A10B25_and(A10B25, A10, B25);
and A9B26_and(A9B26, A9, B26);
and A8B27_and(A8B27, A8, B27);
and A7B28_and(A7B28, A7, B28);
and A6B29_and(A6B29, A6, B29);
and A5B30_and(A5B30, A5, B30);
and A4B31_and(A4B31, A4, B31);

// bit position 35------------------------------------------------------------

wire A31B5, A30B6, A29B7, A28B8, A27B9, A26B10, A25B11, A24B12, A23B13, A22B14, A21B15, A20B16, A19B17, A18B18, A17B19, A16B20, A15B21, A14B22, A13B23, A12B24, A11B25, A10B26, A9B27, A8B28, A7B29, A6B30, A5B31;

and A31B5_and(A31B5, A31, B5);
and A30B6_and(A30B6, A30, B6);
and A29B7_and(A29B7, A29, B7);
and A28B8_and(A28B8, A28, B8);
and A27B9_and(A27B9, A27, B9);
and A26B10_and(A26B10, A26, B10);
and A25B11_and(A25B11, A25, B11);
and A24B12_and(A24B12, A24, B12);
and A23B13_and(A23B13, A23, B13);
and A22B14_and(A22B14, A22, B14);
and A21B15_and(A21B15, A21, B15);
and A20B16_and(A20B16, A20, B16);
and A19B17_and(A19B17, A19, B17);
and A18B18_and(A18B18, A18, B18);
and A17B19_and(A17B19, A17, B19);
and A16B20_and(A16B20, A16, B20);
and A15B21_and(A15B21, A15, B21);
and A14B22_and(A14B22, A14, B22);
and A13B23_and(A13B23, A13, B23);
and A12B24_and(A12B24, A12, B24);
and A11B25_and(A11B25, A11, B25);
and A10B26_and(A10B26, A10, B26);
and A9B27_and(A9B27, A9, B27);
and A8B28_and(A8B28, A8, B28);
and A7B29_and(A7B29, A7, B29);
and A6B30_and(A6B30, A6, B30);
and A5B31_and(A5B31, A5, B31);

// bit position 36------------------------------------------------------------

wire A31B6, A30B7, A29B8, A28B9, A27B10, A26B11, A25B12, A24B13, A23B14, A22B15, A21B16, A20B17, A19B18, A18B19, A17B20, A16B21, A15B22, A14B23, A13B24, A12B25, A11B26, A10B27, A9B28, A8B29, A7B30, A6B31;

and A31B6_and(A31B6, A31, B6);
and A30B7_and(A30B7, A30, B7);
and A29B8_and(A29B8, A29, B8);
and A28B9_and(A28B9, A28, B9);
and A27B10_and(A27B10, A27, B10);
and A26B11_and(A26B11, A26, B11);
and A25B12_and(A25B12, A25, B12);
and A24B13_and(A24B13, A24, B13);
and A23B14_and(A23B14, A23, B14);
and A22B15_and(A22B15, A22, B15);
and A21B16_and(A21B16, A21, B16);
and A20B17_and(A20B17, A20, B17);
and A19B18_and(A19B18, A19, B18);
and A18B19_and(A18B19, A18, B19);
and A17B20_and(A17B20, A17, B20);
and A16B21_and(A16B21, A16, B21);
and A15B22_and(A15B22, A15, B22);
and A14B23_and(A14B23, A14, B23);
and A13B24_and(A13B24, A13, B24);
and A12B25_and(A12B25, A12, B25);
and A11B26_and(A11B26, A11, B26);
and A10B27_and(A10B27, A10, B27);
and A9B28_and(A9B28, A9, B28);
and A8B29_and(A8B29, A8, B29);
and A7B30_and(A7B30, A7, B30);
and A6B31_and(A6B31, A6, B31);

// bit position 37------------------------------------------------------------

wire A31B7, A30B8, A29B9, A28B10, A27B11, A26B12, A25B13, A24B14, A23B15, A22B16, A21B17, A20B18, A19B19, A18B20, A17B21, A16B22, A15B23, A14B24, A13B25, A12B26, A11B27, A10B28, A9B29, A8B30, A7B31;

and A31B7_and(A31B7, A31, B7);
and A30B8_and(A30B8, A30, B8);
and A29B9_and(A29B9, A29, B9);
and A28B10_and(A28B10, A28, B10);
and A27B11_and(A27B11, A27, B11);
and A26B12_and(A26B12, A26, B12);
and A25B13_and(A25B13, A25, B13);
and A24B14_and(A24B14, A24, B14);
and A23B15_and(A23B15, A23, B15);
and A22B16_and(A22B16, A22, B16);
and A21B17_and(A21B17, A21, B17);
and A20B18_and(A20B18, A20, B18);
and A19B19_and(A19B19, A19, B19);
and A18B20_and(A18B20, A18, B20);
and A17B21_and(A17B21, A17, B21);
and A16B22_and(A16B22, A16, B22);
and A15B23_and(A15B23, A15, B23);
and A14B24_and(A14B24, A14, B24);
and A13B25_and(A13B25, A13, B25);
and A12B26_and(A12B26, A12, B26);
and A11B27_and(A11B27, A11, B27);
and A10B28_and(A10B28, A10, B28);
and A9B29_and(A9B29, A9, B29);
and A8B30_and(A8B30, A8, B30);
and A7B31_and(A7B31, A7, B31);

// bit position 38------------------------------------------------------------

wire A31B8, A30B9, A29B10, A28B11, A27B12, A26B13, A25B14, A24B15, A23B16, A22B17, A21B18, A20B19, A19B20, A18B21, A17B22, A16B23, A15B24, A14B25, A13B26, A12B27, A11B28, A10B29, A9B30, A8B31;

and A31B8_and(A31B8, A31, B8);
and A30B9_and(A30B9, A30, B9);
and A29B10_and(A29B10, A29, B10);
and A28B11_and(A28B11, A28, B11);
and A27B12_and(A27B12, A27, B12);
and A26B13_and(A26B13, A26, B13);
and A25B14_and(A25B14, A25, B14);
and A24B15_and(A24B15, A24, B15);
and A23B16_and(A23B16, A23, B16);
and A22B17_and(A22B17, A22, B17);
and A21B18_and(A21B18, A21, B18);
and A20B19_and(A20B19, A20, B19);
and A19B20_and(A19B20, A19, B20);
and A18B21_and(A18B21, A18, B21);
and A17B22_and(A17B22, A17, B22);
and A16B23_and(A16B23, A16, B23);
and A15B24_and(A15B24, A15, B24);
and A14B25_and(A14B25, A14, B25);
and A13B26_and(A13B26, A13, B26);
and A12B27_and(A12B27, A12, B27);
and A11B28_and(A11B28, A11, B28);
and A10B29_and(A10B29, A10, B29);
and A9B30_and(A9B30, A9, B30);
and A8B31_and(A8B31, A8, B31);

// bit position 39------------------------------------------------------------

wire A31B9, A30B10, A29B11, A28B12, A27B13, A26B14, A25B15, A24B16, A23B17, A22B18, A21B19, A20B20, A19B21, A18B22, A17B23, A16B24, A15B25, A14B26, A13B27, A12B28, A11B29, A10B30, A9B31;

and A31B9_and(A31B9, A31, B9);
and A30B10_and(A30B10, A30, B10);
and A29B11_and(A29B11, A29, B11);
and A28B12_and(A28B12, A28, B12);
and A27B13_and(A27B13, A27, B13);
and A26B14_and(A26B14, A26, B14);
and A25B15_and(A25B15, A25, B15);
and A24B16_and(A24B16, A24, B16);
and A23B17_and(A23B17, A23, B17);
and A22B18_and(A22B18, A22, B18);
and A21B19_and(A21B19, A21, B19);
and A20B20_and(A20B20, A20, B20);
and A19B21_and(A19B21, A19, B21);
and A18B22_and(A18B22, A18, B22);
and A17B23_and(A17B23, A17, B23);
and A16B24_and(A16B24, A16, B24);
and A15B25_and(A15B25, A15, B25);
and A14B26_and(A14B26, A14, B26);
and A13B27_and(A13B27, A13, B27);
and A12B28_and(A12B28, A12, B28);
and A11B29_and(A11B29, A11, B29);
and A10B30_and(A10B30, A10, B30);
and A9B31_and(A9B31, A9, B31);

// bit position 40------------------------------------------------------------

wire A31B10, A30B11, A29B12, A28B13, A27B14, A26B15, A25B16, A24B17, A23B18, A22B19, A21B20, A20B21, A19B22, A18B23, A17B24, A16B25, A15B26, A14B27, A13B28, A12B29, A11B30, A10B31;

and A31B10_and(A31B10, A31, B10);
and A30B11_and(A30B11, A30, B11);
and A29B12_and(A29B12, A29, B12);
and A28B13_and(A28B13, A28, B13);
and A27B14_and(A27B14, A27, B14);
and A26B15_and(A26B15, A26, B15);
and A25B16_and(A25B16, A25, B16);
and A24B17_and(A24B17, A24, B17);
and A23B18_and(A23B18, A23, B18);
and A22B19_and(A22B19, A22, B19);
and A21B20_and(A21B20, A21, B20);
and A20B21_and(A20B21, A20, B21);
and A19B22_and(A19B22, A19, B22);
and A18B23_and(A18B23, A18, B23);
and A17B24_and(A17B24, A17, B24);
and A16B25_and(A16B25, A16, B25);
and A15B26_and(A15B26, A15, B26);
and A14B27_and(A14B27, A14, B27);
and A13B28_and(A13B28, A13, B28);
and A12B29_and(A12B29, A12, B29);
and A11B30_and(A11B30, A11, B30);
and A10B31_and(A10B31, A10, B31);

// bit position 41------------------------------------------------------------

wire A31B11, A30B12, A29B13, A28B14, A27B15, A26B16, A25B17, A24B18, A23B19, A22B20, A21B21, A20B22, A19B23, A18B24, A17B25, A16B26, A15B27, A14B28, A13B29, A12B30, A11B31;

and A31B11_and(A31B11, A31, B11);
and A30B12_and(A30B12, A30, B12);
and A29B13_and(A29B13, A29, B13);
and A28B14_and(A28B14, A28, B14);
and A27B15_and(A27B15, A27, B15);
and A26B16_and(A26B16, A26, B16);
and A25B17_and(A25B17, A25, B17);
and A24B18_and(A24B18, A24, B18);
and A23B19_and(A23B19, A23, B19);
and A22B20_and(A22B20, A22, B20);
and A21B21_and(A21B21, A21, B21);
and A20B22_and(A20B22, A20, B22);
and A19B23_and(A19B23, A19, B23);
and A18B24_and(A18B24, A18, B24);
and A17B25_and(A17B25, A17, B25);
and A16B26_and(A16B26, A16, B26);
and A15B27_and(A15B27, A15, B27);
and A14B28_and(A14B28, A14, B28);
and A13B29_and(A13B29, A13, B29);
and A12B30_and(A12B30, A12, B30);
and A11B31_and(A11B31, A11, B31);

// bit position 42------------------------------------------------------------

wire A31B12, A30B13, A29B14, A28B15, A27B16, A26B17, A25B18, A24B19, A23B20, A22B21, A21B22, A20B23, A19B24, A18B25, A17B26, A16B27, A15B28, A14B29, A13B30, A12B31;

and A31B12_and(A31B12, A31, B12);
and A30B13_and(A30B13, A30, B13);
and A29B14_and(A29B14, A29, B14);
and A28B15_and(A28B15, A28, B15);
and A27B16_and(A27B16, A27, B16);
and A26B17_and(A26B17, A26, B17);
and A25B18_and(A25B18, A25, B18);
and A24B19_and(A24B19, A24, B19);
and A23B20_and(A23B20, A23, B20);
and A22B21_and(A22B21, A22, B21);
and A21B22_and(A21B22, A21, B22);
and A20B23_and(A20B23, A20, B23);
and A19B24_and(A19B24, A19, B24);
and A18B25_and(A18B25, A18, B25);
and A17B26_and(A17B26, A17, B26);
and A16B27_and(A16B27, A16, B27);
and A15B28_and(A15B28, A15, B28);
and A14B29_and(A14B29, A14, B29);
and A13B30_and(A13B30, A13, B30);
and A12B31_and(A12B31, A12, B31);

// bit position 43------------------------------------------------------------

wire A31B13, A30B14, A29B15, A28B16, A27B17, A26B18, A25B19, A24B20, A23B21, A22B22, A21B23, A20B24, A19B25, A18B26, A17B27, A16B28, A15B29, A14B30, A13B31;

and A31B13_and(A31B13, A31, B13);
and A30B14_and(A30B14, A30, B14);
and A29B15_and(A29B15, A29, B15);
and A28B16_and(A28B16, A28, B16);
and A27B17_and(A27B17, A27, B17);
and A26B18_and(A26B18, A26, B18);
and A25B19_and(A25B19, A25, B19);
and A24B20_and(A24B20, A24, B20);
and A23B21_and(A23B21, A23, B21);
and A22B22_and(A22B22, A22, B22);
and A21B23_and(A21B23, A21, B23);
and A20B24_and(A20B24, A20, B24);
and A19B25_and(A19B25, A19, B25);
and A18B26_and(A18B26, A18, B26);
and A17B27_and(A17B27, A17, B27);
and A16B28_and(A16B28, A16, B28);
and A15B29_and(A15B29, A15, B29);
and A14B30_and(A14B30, A14, B30);
and A13B31_and(A13B31, A13, B31);

// bit position 44------------------------------------------------------------

wire A31B14, A30B15, A29B16, A28B17, A27B18, A26B19, A25B20, A24B21, A23B22, A22B23, A21B24, A20B25, A19B26, A18B27, A17B28, A16B29, A15B30, A14B31;

and A31B14_and(A31B14, A31, B14);
and A30B15_and(A30B15, A30, B15);
and A29B16_and(A29B16, A29, B16);
and A28B17_and(A28B17, A28, B17);
and A27B18_and(A27B18, A27, B18);
and A26B19_and(A26B19, A26, B19);
and A25B20_and(A25B20, A25, B20);
and A24B21_and(A24B21, A24, B21);
and A23B22_and(A23B22, A23, B22);
and A22B23_and(A22B23, A22, B23);
and A21B24_and(A21B24, A21, B24);
and A20B25_and(A20B25, A20, B25);
and A19B26_and(A19B26, A19, B26);
and A18B27_and(A18B27, A18, B27);
and A17B28_and(A17B28, A17, B28);
and A16B29_and(A16B29, A16, B29);
and A15B30_and(A15B30, A15, B30);
and A14B31_and(A14B31, A14, B31);

// bit position 45------------------------------------------------------------

wire A31B15, A30B16, A29B17, A28B18, A27B19, A26B20, A25B21, A24B22, A23B23, A22B24, A21B25, A20B26, A19B27, A18B28, A17B29, A16B30, A15B31;

and A31B15_and(A31B15, A31, B15);
and A30B16_and(A30B16, A30, B16);
and A29B17_and(A29B17, A29, B17);
and A28B18_and(A28B18, A28, B18);
and A27B19_and(A27B19, A27, B19);
and A26B20_and(A26B20, A26, B20);
and A25B21_and(A25B21, A25, B21);
and A24B22_and(A24B22, A24, B22);
and A23B23_and(A23B23, A23, B23);
and A22B24_and(A22B24, A22, B24);
and A21B25_and(A21B25, A21, B25);
and A20B26_and(A20B26, A20, B26);
and A19B27_and(A19B27, A19, B27);
and A18B28_and(A18B28, A18, B28);
and A17B29_and(A17B29, A17, B29);
and A16B30_and(A16B30, A16, B30);
and A15B31_and(A15B31, A15, B31);

// bit position 46------------------------------------------------------------

wire A31B16, A30B17, A29B18, A28B19, A27B20, A26B21, A25B22, A24B23, A23B24, A22B25, A21B26, A20B27, A19B28, A18B29, A17B30, A16B31;

and A31B16_and(A31B16, A31, B16);
and A30B17_and(A30B17, A30, B17);
and A29B18_and(A29B18, A29, B18);
and A28B19_and(A28B19, A28, B19);
and A27B20_and(A27B20, A27, B20);
and A26B21_and(A26B21, A26, B21);
and A25B22_and(A25B22, A25, B22);
and A24B23_and(A24B23, A24, B23);
and A23B24_and(A23B24, A23, B24);
and A22B25_and(A22B25, A22, B25);
and A21B26_and(A21B26, A21, B26);
and A20B27_and(A20B27, A20, B27);
and A19B28_and(A19B28, A19, B28);
and A18B29_and(A18B29, A18, B29);
and A17B30_and(A17B30, A17, B30);
and A16B31_and(A16B31, A16, B31);

// bit position 47------------------------------------------------------------

wire A31B17, A30B18, A29B19, A28B20, A27B21, A26B22, A25B23, A24B24, A23B25, A22B26, A21B27, A20B28, A19B29, A18B30, A17B31;

and A31B17_and(A31B17, A31, B17);
and A30B18_and(A30B18, A30, B18);
and A29B19_and(A29B19, A29, B19);
and A28B20_and(A28B20, A28, B20);
and A27B21_and(A27B21, A27, B21);
and A26B22_and(A26B22, A26, B22);
and A25B23_and(A25B23, A25, B23);
and A24B24_and(A24B24, A24, B24);
and A23B25_and(A23B25, A23, B25);
and A22B26_and(A22B26, A22, B26);
and A21B27_and(A21B27, A21, B27);
and A20B28_and(A20B28, A20, B28);
and A19B29_and(A19B29, A19, B29);
and A18B30_and(A18B30, A18, B30);
and A17B31_and(A17B31, A17, B31);

// bit position 48------------------------------------------------------------

wire A31B18, A30B19, A29B20, A28B21, A27B22, A26B23, A25B24, A24B25, A23B26, A22B27, A21B28, A20B29, A19B30, A18B31;

and A31B18_and(A31B18, A31, B18);
and A30B19_and(A30B19, A30, B19);
and A29B20_and(A29B20, A29, B20);
and A28B21_and(A28B21, A28, B21);
and A27B22_and(A27B22, A27, B22);
and A26B23_and(A26B23, A26, B23);
and A25B24_and(A25B24, A25, B24);
and A24B25_and(A24B25, A24, B25);
and A23B26_and(A23B26, A23, B26);
and A22B27_and(A22B27, A22, B27);
and A21B28_and(A21B28, A21, B28);
and A20B29_and(A20B29, A20, B29);
and A19B30_and(A19B30, A19, B30);
and A18B31_and(A18B31, A18, B31);

// bit position 49------------------------------------------------------------

wire A31B19, A30B20, A29B21, A28B22, A27B23, A26B24, A25B25, A24B26, A23B27, A22B28, A21B29, A20B30, A19B31;

and A31B19_and(A31B19, A31, B19);
and A30B20_and(A30B20, A30, B20);
and A29B21_and(A29B21, A29, B21);
and A28B22_and(A28B22, A28, B22);
and A27B23_and(A27B23, A27, B23);
and A26B24_and(A26B24, A26, B24);
and A25B25_and(A25B25, A25, B25);
and A24B26_and(A24B26, A24, B26);
and A23B27_and(A23B27, A23, B27);
and A22B28_and(A22B28, A22, B28);
and A21B29_and(A21B29, A21, B29);
and A20B30_and(A20B30, A20, B30);
and A19B31_and(A19B31, A19, B31);

// bit position 50------------------------------------------------------------

wire A31B20, A30B21, A29B22, A28B23, A27B24, A26B25, A25B26, A24B27, A23B28, A22B29, A21B30, A20B31;

and A31B20_and(A31B20, A31, B20);
and A30B21_and(A30B21, A30, B21);
and A29B22_and(A29B22, A29, B22);
and A28B23_and(A28B23, A28, B23);
and A27B24_and(A27B24, A27, B24);
and A26B25_and(A26B25, A26, B25);
and A25B26_and(A25B26, A25, B26);
and A24B27_and(A24B27, A24, B27);
and A23B28_and(A23B28, A23, B28);
and A22B29_and(A22B29, A22, B29);
and A21B30_and(A21B30, A21, B30);
and A20B31_and(A20B31, A20, B31);

// bit position 51------------------------------------------------------------

wire A31B21, A30B22, A29B23, A28B24, A27B25, A26B26, A25B27, A24B28, A23B29, A22B30, A21B31;

and A31B21_and(A31B21, A31, B21);
and A30B22_and(A30B22, A30, B22);
and A29B23_and(A29B23, A29, B23);
and A28B24_and(A28B24, A28, B24);
and A27B25_and(A27B25, A27, B25);
and A26B26_and(A26B26, A26, B26);
and A25B27_and(A25B27, A25, B27);
and A24B28_and(A24B28, A24, B28);
and A23B29_and(A23B29, A23, B29);
and A22B30_and(A22B30, A22, B30);
and A21B31_and(A21B31, A21, B31);

// bit position 52------------------------------------------------------------

wire A31B22, A30B23, A29B24, A28B25, A27B26, A26B27, A25B28, A24B29, A23B30, A22B31;

and A31B22_and(A31B22, A31, B22);
and A30B23_and(A30B23, A30, B23);
and A29B24_and(A29B24, A29, B24);
and A28B25_and(A28B25, A28, B25);
and A27B26_and(A27B26, A27, B26);
and A26B27_and(A26B27, A26, B27);
and A25B28_and(A25B28, A25, B28);
and A24B29_and(A24B29, A24, B29);
and A23B30_and(A23B30, A23, B30);
and A22B31_and(A22B31, A22, B31);

// bit position 53------------------------------------------------------------

wire A31B23, A30B24, A29B25, A28B26, A27B27, A26B28, A25B29, A24B30, A23B31;

and A31B23_and(A31B23, A31, B23);
and A30B24_and(A30B24, A30, B24);
and A29B25_and(A29B25, A29, B25);
and A28B26_and(A28B26, A28, B26);
and A27B27_and(A27B27, A27, B27);
and A26B28_and(A26B28, A26, B28);
and A25B29_and(A25B29, A25, B29);
and A24B30_and(A24B30, A24, B30);
and A23B31_and(A23B31, A23, B31);

// bit position 54------------------------------------------------------------

wire A31B24, A30B25, A29B26, A28B27, A27B28, A26B29, A25B30, A24B31;

and A31B24_and(A31B24, A31, B24);
and A30B25_and(A30B25, A30, B25);
and A29B26_and(A29B26, A29, B26);
and A28B27_and(A28B27, A28, B27);
and A27B28_and(A27B28, A27, B28);
and A26B29_and(A26B29, A26, B29);
and A25B30_and(A25B30, A25, B30);
and A24B31_and(A24B31, A24, B31);

// bit position 55------------------------------------------------------------

wire A31B25, A30B26, A29B27, A28B28, A27B29, A26B30, A25B31;

and A31B25_and(A31B25, A31, B25);
and A30B26_and(A30B26, A30, B26);
and A29B27_and(A29B27, A29, B27);
and A28B28_and(A28B28, A28, B28);
and A27B29_and(A27B29, A27, B29);
and A26B30_and(A26B30, A26, B30);
and A25B31_and(A25B31, A25, B31);

// bit position 56------------------------------------------------------------

wire A31B26, A30B27, A29B28, A28B29, A27B30, A26B31;

and A31B26_and(A31B26, A31, B26);
and A30B27_and(A30B27, A30, B27);
and A29B28_and(A29B28, A29, B28);
and A28B29_and(A28B29, A28, B29);
and A27B30_and(A27B30, A27, B30);
and A26B31_and(A26B31, A26, B31);

// bit position 57------------------------------------------------------------

wire A31B27, A30B28, A29B29, A28B30, A27B31;

and A31B27_and(A31B27, A31, B27);
and A30B28_and(A30B28, A30, B28);
and A29B29_and(A29B29, A29, B29);
and A28B30_and(A28B30, A28, B30);
and A27B31_and(A27B31, A27, B31);

// bit position 58------------------------------------------------------------

wire A31B28, A30B29, A29B30, A28B31;

and A31B28_and(A31B28, A31, B28);
and A30B29_and(A30B29, A30, B29);
and A29B30_and(A29B30, A29, B30);
and A28B31_and(A28B31, A28, B31);

// bit position 59------------------------------------------------------------

wire A31B29, A30B30, A29B31;

and A31B29_and(A31B29, A31, B29);
and A30B30_and(A30B30, A30, B30);
and A29B31_and(A29B31, A29, B31);

// bit position 60------------------------------------------------------------

wire A31B30, A30B31;

and A31B30_and(A31B30, A31, B30);
and A30B31_and(A30B31, A30, B31);

// bit position 61------------------------------------------------------------

wire A31B31;

and A31B31_and(A31B31, A31, B31);

// bit position 62------------------------------------------------------------

wire sum_2_0_0, cout_2_0_0;

half_adder ha_2_0_0(sum_2_0_0, cout_2_0_0, A2B0, A1B1);

wire sum_3_0_0, cout_3_0_0;

full_adder fa_3_0_0(sum_3_0_0, cout_3_0_0, A3B0, A2B1, A1B2);

wire sum_4_0_0, cout_4_0_0;

full_adder fa_4_0_0(sum_4_0_0, cout_4_0_0, A4B0, A3B1, A2B2);

wire sum_4_1_0, cout_4_1_0;

half_adder ha_4_1_0(sum_4_1_0, cout_4_1_0, A1B3, A0B4);

wire sum_5_0_0, cout_5_0_0;

full_adder fa_5_0_0(sum_5_0_0, cout_5_0_0, A5B0, A4B1, A3B2);

wire sum_5_1_0, cout_5_1_0;

full_adder fa_5_1_0(sum_5_1_0, cout_5_1_0, A2B3, A1B4, A0B5);

wire sum_6_0_0, cout_6_0_0;

full_adder fa_6_0_0(sum_6_0_0, cout_6_0_0, A6B0, A5B1, A4B2);

wire sum_6_1_0, cout_6_1_0;

full_adder fa_6_1_0(sum_6_1_0, cout_6_1_0, A3B3, A2B4, A1B5);

wire sum_7_0_0, cout_7_0_0;

full_adder fa_7_0_0(sum_7_0_0, cout_7_0_0, A7B0, A6B1, A5B2);

wire sum_7_1_0, cout_7_1_0;

full_adder fa_7_1_0(sum_7_1_0, cout_7_1_0, A4B3, A3B4, A2B5);

wire sum_7_2_0, cout_7_2_0;

half_adder ha_7_2_0(sum_7_2_0, cout_7_2_0, A1B6, A0B7);

wire sum_8_0_0, cout_8_0_0;

full_adder fa_8_0_0(sum_8_0_0, cout_8_0_0, A8B0, A7B1, A6B2);

wire sum_8_1_0, cout_8_1_0;

full_adder fa_8_1_0(sum_8_1_0, cout_8_1_0, A5B3, A4B4, A3B5);

wire sum_8_2_0, cout_8_2_0;

full_adder fa_8_2_0(sum_8_2_0, cout_8_2_0, A2B6, A1B7, A0B8);

wire sum_9_0_0, cout_9_0_0;

full_adder fa_9_0_0(sum_9_0_0, cout_9_0_0, A9B0, A8B1, A7B2);

wire sum_9_1_0, cout_9_1_0;

full_adder fa_9_1_0(sum_9_1_0, cout_9_1_0, A6B3, A5B4, A4B5);

wire sum_9_2_0, cout_9_2_0;

full_adder fa_9_2_0(sum_9_2_0, cout_9_2_0, A3B6, A2B7, A1B8);

wire sum_10_0_0, cout_10_0_0;

full_adder fa_10_0_0(sum_10_0_0, cout_10_0_0, A10B0, A9B1, A8B2);

wire sum_10_1_0, cout_10_1_0;

full_adder fa_10_1_0(sum_10_1_0, cout_10_1_0, A7B3, A6B4, A5B5);

wire sum_10_2_0, cout_10_2_0;

full_adder fa_10_2_0(sum_10_2_0, cout_10_2_0, A4B6, A3B7, A2B8);

wire sum_10_3_0, cout_10_3_0;

half_adder ha_10_3_0(sum_10_3_0, cout_10_3_0, A1B9, A0B10);

wire sum_11_0_0, cout_11_0_0;

full_adder fa_11_0_0(sum_11_0_0, cout_11_0_0, A11B0, A10B1, A9B2);

wire sum_11_1_0, cout_11_1_0;

full_adder fa_11_1_0(sum_11_1_0, cout_11_1_0, A8B3, A7B4, A6B5);

wire sum_11_2_0, cout_11_2_0;

full_adder fa_11_2_0(sum_11_2_0, cout_11_2_0, A5B6, A4B7, A3B8);

wire sum_11_3_0, cout_11_3_0;

full_adder fa_11_3_0(sum_11_3_0, cout_11_3_0, A2B9, A1B10, A0B11);

wire sum_12_0_0, cout_12_0_0;

full_adder fa_12_0_0(sum_12_0_0, cout_12_0_0, A12B0, A11B1, A10B2);

wire sum_12_1_0, cout_12_1_0;

full_adder fa_12_1_0(sum_12_1_0, cout_12_1_0, A9B3, A8B4, A7B5);

wire sum_12_2_0, cout_12_2_0;

full_adder fa_12_2_0(sum_12_2_0, cout_12_2_0, A6B6, A5B7, A4B8);

wire sum_12_3_0, cout_12_3_0;

full_adder fa_12_3_0(sum_12_3_0, cout_12_3_0, A3B9, A2B10, A1B11);

wire sum_13_0_0, cout_13_0_0;

full_adder fa_13_0_0(sum_13_0_0, cout_13_0_0, A13B0, A12B1, A11B2);

wire sum_13_1_0, cout_13_1_0;

full_adder fa_13_1_0(sum_13_1_0, cout_13_1_0, A10B3, A9B4, A8B5);

wire sum_13_2_0, cout_13_2_0;

full_adder fa_13_2_0(sum_13_2_0, cout_13_2_0, A7B6, A6B7, A5B8);

wire sum_13_3_0, cout_13_3_0;

full_adder fa_13_3_0(sum_13_3_0, cout_13_3_0, A4B9, A3B10, A2B11);

wire sum_13_4_0, cout_13_4_0;

half_adder ha_13_4_0(sum_13_4_0, cout_13_4_0, A1B12, A0B13);

wire sum_14_0_0, cout_14_0_0;

full_adder fa_14_0_0(sum_14_0_0, cout_14_0_0, A14B0, A13B1, A12B2);

wire sum_14_1_0, cout_14_1_0;

full_adder fa_14_1_0(sum_14_1_0, cout_14_1_0, A11B3, A10B4, A9B5);

wire sum_14_2_0, cout_14_2_0;

full_adder fa_14_2_0(sum_14_2_0, cout_14_2_0, A8B6, A7B7, A6B8);

wire sum_14_3_0, cout_14_3_0;

full_adder fa_14_3_0(sum_14_3_0, cout_14_3_0, A5B9, A4B10, A3B11);

wire sum_14_4_0, cout_14_4_0;

full_adder fa_14_4_0(sum_14_4_0, cout_14_4_0, A2B12, A1B13, A0B14);

wire sum_15_0_0, cout_15_0_0;

full_adder fa_15_0_0(sum_15_0_0, cout_15_0_0, A15B0, A14B1, A13B2);

wire sum_15_1_0, cout_15_1_0;

full_adder fa_15_1_0(sum_15_1_0, cout_15_1_0, A12B3, A11B4, A10B5);

wire sum_15_2_0, cout_15_2_0;

full_adder fa_15_2_0(sum_15_2_0, cout_15_2_0, A9B6, A8B7, A7B8);

wire sum_15_3_0, cout_15_3_0;

full_adder fa_15_3_0(sum_15_3_0, cout_15_3_0, A6B9, A5B10, A4B11);

wire sum_15_4_0, cout_15_4_0;

full_adder fa_15_4_0(sum_15_4_0, cout_15_4_0, A3B12, A2B13, A1B14);

wire sum_16_0_0, cout_16_0_0;

full_adder fa_16_0_0(sum_16_0_0, cout_16_0_0, A16B0, A15B1, A14B2);

wire sum_16_1_0, cout_16_1_0;

full_adder fa_16_1_0(sum_16_1_0, cout_16_1_0, A13B3, A12B4, A11B5);

wire sum_16_2_0, cout_16_2_0;

full_adder fa_16_2_0(sum_16_2_0, cout_16_2_0, A10B6, A9B7, A8B8);

wire sum_16_3_0, cout_16_3_0;

full_adder fa_16_3_0(sum_16_3_0, cout_16_3_0, A7B9, A6B10, A5B11);

wire sum_16_4_0, cout_16_4_0;

full_adder fa_16_4_0(sum_16_4_0, cout_16_4_0, A4B12, A3B13, A2B14);

wire sum_16_5_0, cout_16_5_0;

half_adder ha_16_5_0(sum_16_5_0, cout_16_5_0, A1B15, A0B16);

wire sum_17_0_0, cout_17_0_0;

full_adder fa_17_0_0(sum_17_0_0, cout_17_0_0, A17B0, A16B1, A15B2);

wire sum_17_1_0, cout_17_1_0;

full_adder fa_17_1_0(sum_17_1_0, cout_17_1_0, A14B3, A13B4, A12B5);

wire sum_17_2_0, cout_17_2_0;

full_adder fa_17_2_0(sum_17_2_0, cout_17_2_0, A11B6, A10B7, A9B8);

wire sum_17_3_0, cout_17_3_0;

full_adder fa_17_3_0(sum_17_3_0, cout_17_3_0, A8B9, A7B10, A6B11);

wire sum_17_4_0, cout_17_4_0;

full_adder fa_17_4_0(sum_17_4_0, cout_17_4_0, A5B12, A4B13, A3B14);

wire sum_17_5_0, cout_17_5_0;

full_adder fa_17_5_0(sum_17_5_0, cout_17_5_0, A2B15, A1B16, A0B17);

wire sum_18_0_0, cout_18_0_0;

full_adder fa_18_0_0(sum_18_0_0, cout_18_0_0, A18B0, A17B1, A16B2);

wire sum_18_1_0, cout_18_1_0;

full_adder fa_18_1_0(sum_18_1_0, cout_18_1_0, A15B3, A14B4, A13B5);

wire sum_18_2_0, cout_18_2_0;

full_adder fa_18_2_0(sum_18_2_0, cout_18_2_0, A12B6, A11B7, A10B8);

wire sum_18_3_0, cout_18_3_0;

full_adder fa_18_3_0(sum_18_3_0, cout_18_3_0, A9B9, A8B10, A7B11);

wire sum_18_4_0, cout_18_4_0;

full_adder fa_18_4_0(sum_18_4_0, cout_18_4_0, A6B12, A5B13, A4B14);

wire sum_18_5_0, cout_18_5_0;

full_adder fa_18_5_0(sum_18_5_0, cout_18_5_0, A3B15, A2B16, A1B17);

wire sum_19_0_0, cout_19_0_0;

full_adder fa_19_0_0(sum_19_0_0, cout_19_0_0, A19B0, A18B1, A17B2);

wire sum_19_1_0, cout_19_1_0;

full_adder fa_19_1_0(sum_19_1_0, cout_19_1_0, A16B3, A15B4, A14B5);

wire sum_19_2_0, cout_19_2_0;

full_adder fa_19_2_0(sum_19_2_0, cout_19_2_0, A13B6, A12B7, A11B8);

wire sum_19_3_0, cout_19_3_0;

full_adder fa_19_3_0(sum_19_3_0, cout_19_3_0, A10B9, A9B10, A8B11);

wire sum_19_4_0, cout_19_4_0;

full_adder fa_19_4_0(sum_19_4_0, cout_19_4_0, A7B12, A6B13, A5B14);

wire sum_19_5_0, cout_19_5_0;

full_adder fa_19_5_0(sum_19_5_0, cout_19_5_0, A4B15, A3B16, A2B17);

wire sum_19_6_0, cout_19_6_0;

half_adder ha_19_6_0(sum_19_6_0, cout_19_6_0, A1B18, A0B19);

wire sum_20_0_0, cout_20_0_0;

full_adder fa_20_0_0(sum_20_0_0, cout_20_0_0, A20B0, A19B1, A18B2);

wire sum_20_1_0, cout_20_1_0;

full_adder fa_20_1_0(sum_20_1_0, cout_20_1_0, A17B3, A16B4, A15B5);

wire sum_20_2_0, cout_20_2_0;

full_adder fa_20_2_0(sum_20_2_0, cout_20_2_0, A14B6, A13B7, A12B8);

wire sum_20_3_0, cout_20_3_0;

full_adder fa_20_3_0(sum_20_3_0, cout_20_3_0, A11B9, A10B10, A9B11);

wire sum_20_4_0, cout_20_4_0;

full_adder fa_20_4_0(sum_20_4_0, cout_20_4_0, A8B12, A7B13, A6B14);

wire sum_20_5_0, cout_20_5_0;

full_adder fa_20_5_0(sum_20_5_0, cout_20_5_0, A5B15, A4B16, A3B17);

wire sum_20_6_0, cout_20_6_0;

full_adder fa_20_6_0(sum_20_6_0, cout_20_6_0, A2B18, A1B19, A0B20);

wire sum_21_0_0, cout_21_0_0;

full_adder fa_21_0_0(sum_21_0_0, cout_21_0_0, A21B0, A20B1, A19B2);

wire sum_21_1_0, cout_21_1_0;

full_adder fa_21_1_0(sum_21_1_0, cout_21_1_0, A18B3, A17B4, A16B5);

wire sum_21_2_0, cout_21_2_0;

full_adder fa_21_2_0(sum_21_2_0, cout_21_2_0, A15B6, A14B7, A13B8);

wire sum_21_3_0, cout_21_3_0;

full_adder fa_21_3_0(sum_21_3_0, cout_21_3_0, A12B9, A11B10, A10B11);

wire sum_21_4_0, cout_21_4_0;

full_adder fa_21_4_0(sum_21_4_0, cout_21_4_0, A9B12, A8B13, A7B14);

wire sum_21_5_0, cout_21_5_0;

full_adder fa_21_5_0(sum_21_5_0, cout_21_5_0, A6B15, A5B16, A4B17);

wire sum_21_6_0, cout_21_6_0;

full_adder fa_21_6_0(sum_21_6_0, cout_21_6_0, A3B18, A2B19, A1B20);

wire sum_22_0_0, cout_22_0_0;

full_adder fa_22_0_0(sum_22_0_0, cout_22_0_0, A22B0, A21B1, A20B2);

wire sum_22_1_0, cout_22_1_0;

full_adder fa_22_1_0(sum_22_1_0, cout_22_1_0, A19B3, A18B4, A17B5);

wire sum_22_2_0, cout_22_2_0;

full_adder fa_22_2_0(sum_22_2_0, cout_22_2_0, A16B6, A15B7, A14B8);

wire sum_22_3_0, cout_22_3_0;

full_adder fa_22_3_0(sum_22_3_0, cout_22_3_0, A13B9, A12B10, A11B11);

wire sum_22_4_0, cout_22_4_0;

full_adder fa_22_4_0(sum_22_4_0, cout_22_4_0, A10B12, A9B13, A8B14);

wire sum_22_5_0, cout_22_5_0;

full_adder fa_22_5_0(sum_22_5_0, cout_22_5_0, A7B15, A6B16, A5B17);

wire sum_22_6_0, cout_22_6_0;

full_adder fa_22_6_0(sum_22_6_0, cout_22_6_0, A4B18, A3B19, A2B20);

wire sum_22_7_0, cout_22_7_0;

half_adder ha_22_7_0(sum_22_7_0, cout_22_7_0, A1B21, A0B22);

wire sum_23_0_0, cout_23_0_0;

full_adder fa_23_0_0(sum_23_0_0, cout_23_0_0, A23B0, A22B1, A21B2);

wire sum_23_1_0, cout_23_1_0;

full_adder fa_23_1_0(sum_23_1_0, cout_23_1_0, A20B3, A19B4, A18B5);

wire sum_23_2_0, cout_23_2_0;

full_adder fa_23_2_0(sum_23_2_0, cout_23_2_0, A17B6, A16B7, A15B8);

wire sum_23_3_0, cout_23_3_0;

full_adder fa_23_3_0(sum_23_3_0, cout_23_3_0, A14B9, A13B10, A12B11);

wire sum_23_4_0, cout_23_4_0;

full_adder fa_23_4_0(sum_23_4_0, cout_23_4_0, A11B12, A10B13, A9B14);

wire sum_23_5_0, cout_23_5_0;

full_adder fa_23_5_0(sum_23_5_0, cout_23_5_0, A8B15, A7B16, A6B17);

wire sum_23_6_0, cout_23_6_0;

full_adder fa_23_6_0(sum_23_6_0, cout_23_6_0, A5B18, A4B19, A3B20);

wire sum_23_7_0, cout_23_7_0;

full_adder fa_23_7_0(sum_23_7_0, cout_23_7_0, A2B21, A1B22, A0B23);

wire sum_24_0_0, cout_24_0_0;

full_adder fa_24_0_0(sum_24_0_0, cout_24_0_0, A24B0, A23B1, A22B2);

wire sum_24_1_0, cout_24_1_0;

full_adder fa_24_1_0(sum_24_1_0, cout_24_1_0, A21B3, A20B4, A19B5);

wire sum_24_2_0, cout_24_2_0;

full_adder fa_24_2_0(sum_24_2_0, cout_24_2_0, A18B6, A17B7, A16B8);

wire sum_24_3_0, cout_24_3_0;

full_adder fa_24_3_0(sum_24_3_0, cout_24_3_0, A15B9, A14B10, A13B11);

wire sum_24_4_0, cout_24_4_0;

full_adder fa_24_4_0(sum_24_4_0, cout_24_4_0, A12B12, A11B13, A10B14);

wire sum_24_5_0, cout_24_5_0;

full_adder fa_24_5_0(sum_24_5_0, cout_24_5_0, A9B15, A8B16, A7B17);

wire sum_24_6_0, cout_24_6_0;

full_adder fa_24_6_0(sum_24_6_0, cout_24_6_0, A6B18, A5B19, A4B20);

wire sum_24_7_0, cout_24_7_0;

full_adder fa_24_7_0(sum_24_7_0, cout_24_7_0, A3B21, A2B22, A1B23);

wire sum_25_0_0, cout_25_0_0;

full_adder fa_25_0_0(sum_25_0_0, cout_25_0_0, A25B0, A24B1, A23B2);

wire sum_25_1_0, cout_25_1_0;

full_adder fa_25_1_0(sum_25_1_0, cout_25_1_0, A22B3, A21B4, A20B5);

wire sum_25_2_0, cout_25_2_0;

full_adder fa_25_2_0(sum_25_2_0, cout_25_2_0, A19B6, A18B7, A17B8);

wire sum_25_3_0, cout_25_3_0;

full_adder fa_25_3_0(sum_25_3_0, cout_25_3_0, A16B9, A15B10, A14B11);

wire sum_25_4_0, cout_25_4_0;

full_adder fa_25_4_0(sum_25_4_0, cout_25_4_0, A13B12, A12B13, A11B14);

wire sum_25_5_0, cout_25_5_0;

full_adder fa_25_5_0(sum_25_5_0, cout_25_5_0, A10B15, A9B16, A8B17);

wire sum_25_6_0, cout_25_6_0;

full_adder fa_25_6_0(sum_25_6_0, cout_25_6_0, A7B18, A6B19, A5B20);

wire sum_25_7_0, cout_25_7_0;

full_adder fa_25_7_0(sum_25_7_0, cout_25_7_0, A4B21, A3B22, A2B23);

wire sum_25_8_0, cout_25_8_0;

half_adder ha_25_8_0(sum_25_8_0, cout_25_8_0, A1B24, A0B25);

wire sum_26_0_0, cout_26_0_0;

full_adder fa_26_0_0(sum_26_0_0, cout_26_0_0, A26B0, A25B1, A24B2);

wire sum_26_1_0, cout_26_1_0;

full_adder fa_26_1_0(sum_26_1_0, cout_26_1_0, A23B3, A22B4, A21B5);

wire sum_26_2_0, cout_26_2_0;

full_adder fa_26_2_0(sum_26_2_0, cout_26_2_0, A20B6, A19B7, A18B8);

wire sum_26_3_0, cout_26_3_0;

full_adder fa_26_3_0(sum_26_3_0, cout_26_3_0, A17B9, A16B10, A15B11);

wire sum_26_4_0, cout_26_4_0;

full_adder fa_26_4_0(sum_26_4_0, cout_26_4_0, A14B12, A13B13, A12B14);

wire sum_26_5_0, cout_26_5_0;

full_adder fa_26_5_0(sum_26_5_0, cout_26_5_0, A11B15, A10B16, A9B17);

wire sum_26_6_0, cout_26_6_0;

full_adder fa_26_6_0(sum_26_6_0, cout_26_6_0, A8B18, A7B19, A6B20);

wire sum_26_7_0, cout_26_7_0;

full_adder fa_26_7_0(sum_26_7_0, cout_26_7_0, A5B21, A4B22, A3B23);

wire sum_26_8_0, cout_26_8_0;

full_adder fa_26_8_0(sum_26_8_0, cout_26_8_0, A2B24, A1B25, A0B26);

wire sum_27_0_0, cout_27_0_0;

full_adder fa_27_0_0(sum_27_0_0, cout_27_0_0, A27B0, A26B1, A25B2);

wire sum_27_1_0, cout_27_1_0;

full_adder fa_27_1_0(sum_27_1_0, cout_27_1_0, A24B3, A23B4, A22B5);

wire sum_27_2_0, cout_27_2_0;

full_adder fa_27_2_0(sum_27_2_0, cout_27_2_0, A21B6, A20B7, A19B8);

wire sum_27_3_0, cout_27_3_0;

full_adder fa_27_3_0(sum_27_3_0, cout_27_3_0, A18B9, A17B10, A16B11);

wire sum_27_4_0, cout_27_4_0;

full_adder fa_27_4_0(sum_27_4_0, cout_27_4_0, A15B12, A14B13, A13B14);

wire sum_27_5_0, cout_27_5_0;

full_adder fa_27_5_0(sum_27_5_0, cout_27_5_0, A12B15, A11B16, A10B17);

wire sum_27_6_0, cout_27_6_0;

full_adder fa_27_6_0(sum_27_6_0, cout_27_6_0, A9B18, A8B19, A7B20);

wire sum_27_7_0, cout_27_7_0;

full_adder fa_27_7_0(sum_27_7_0, cout_27_7_0, A6B21, A5B22, A4B23);

wire sum_27_8_0, cout_27_8_0;

full_adder fa_27_8_0(sum_27_8_0, cout_27_8_0, A3B24, A2B25, A1B26);

wire sum_28_0_0, cout_28_0_0;

full_adder fa_28_0_0(sum_28_0_0, cout_28_0_0, A28B0, A27B1, A26B2);

wire sum_28_1_0, cout_28_1_0;

full_adder fa_28_1_0(sum_28_1_0, cout_28_1_0, A25B3, A24B4, A23B5);

wire sum_28_2_0, cout_28_2_0;

full_adder fa_28_2_0(sum_28_2_0, cout_28_2_0, A22B6, A21B7, A20B8);

wire sum_28_3_0, cout_28_3_0;

full_adder fa_28_3_0(sum_28_3_0, cout_28_3_0, A19B9, A18B10, A17B11);

wire sum_28_4_0, cout_28_4_0;

full_adder fa_28_4_0(sum_28_4_0, cout_28_4_0, A16B12, A15B13, A14B14);

wire sum_28_5_0, cout_28_5_0;

full_adder fa_28_5_0(sum_28_5_0, cout_28_5_0, A13B15, A12B16, A11B17);

wire sum_28_6_0, cout_28_6_0;

full_adder fa_28_6_0(sum_28_6_0, cout_28_6_0, A10B18, A9B19, A8B20);

wire sum_28_7_0, cout_28_7_0;

full_adder fa_28_7_0(sum_28_7_0, cout_28_7_0, A7B21, A6B22, A5B23);

wire sum_28_8_0, cout_28_8_0;

full_adder fa_28_8_0(sum_28_8_0, cout_28_8_0, A4B24, A3B25, A2B26);

wire sum_28_9_0, cout_28_9_0;

half_adder ha_28_9_0(sum_28_9_0, cout_28_9_0, A1B27, A0B28);

wire sum_29_0_0, cout_29_0_0;

full_adder fa_29_0_0(sum_29_0_0, cout_29_0_0, A29B0, A28B1, A27B2);

wire sum_29_1_0, cout_29_1_0;

full_adder fa_29_1_0(sum_29_1_0, cout_29_1_0, A26B3, A25B4, A24B5);

wire sum_29_2_0, cout_29_2_0;

full_adder fa_29_2_0(sum_29_2_0, cout_29_2_0, A23B6, A22B7, A21B8);

wire sum_29_3_0, cout_29_3_0;

full_adder fa_29_3_0(sum_29_3_0, cout_29_3_0, A20B9, A19B10, A18B11);

wire sum_29_4_0, cout_29_4_0;

full_adder fa_29_4_0(sum_29_4_0, cout_29_4_0, A17B12, A16B13, A15B14);

wire sum_29_5_0, cout_29_5_0;

full_adder fa_29_5_0(sum_29_5_0, cout_29_5_0, A14B15, A13B16, A12B17);

wire sum_29_6_0, cout_29_6_0;

full_adder fa_29_6_0(sum_29_6_0, cout_29_6_0, A11B18, A10B19, A9B20);

wire sum_29_7_0, cout_29_7_0;

full_adder fa_29_7_0(sum_29_7_0, cout_29_7_0, A8B21, A7B22, A6B23);

wire sum_29_8_0, cout_29_8_0;

full_adder fa_29_8_0(sum_29_8_0, cout_29_8_0, A5B24, A4B25, A3B26);

wire sum_29_9_0, cout_29_9_0;

full_adder fa_29_9_0(sum_29_9_0, cout_29_9_0, A2B27, A1B28, A0B29);

wire sum_30_0_0, cout_30_0_0;

full_adder fa_30_0_0(sum_30_0_0, cout_30_0_0, A30B0, A29B1, A28B2);

wire sum_30_1_0, cout_30_1_0;

full_adder fa_30_1_0(sum_30_1_0, cout_30_1_0, A27B3, A26B4, A25B5);

wire sum_30_2_0, cout_30_2_0;

full_adder fa_30_2_0(sum_30_2_0, cout_30_2_0, A24B6, A23B7, A22B8);

wire sum_30_3_0, cout_30_3_0;

full_adder fa_30_3_0(sum_30_3_0, cout_30_3_0, A21B9, A20B10, A19B11);

wire sum_30_4_0, cout_30_4_0;

full_adder fa_30_4_0(sum_30_4_0, cout_30_4_0, A18B12, A17B13, A16B14);

wire sum_30_5_0, cout_30_5_0;

full_adder fa_30_5_0(sum_30_5_0, cout_30_5_0, A15B15, A14B16, A13B17);

wire sum_30_6_0, cout_30_6_0;

full_adder fa_30_6_0(sum_30_6_0, cout_30_6_0, A12B18, A11B19, A10B20);

wire sum_30_7_0, cout_30_7_0;

full_adder fa_30_7_0(sum_30_7_0, cout_30_7_0, A9B21, A8B22, A7B23);

wire sum_30_8_0, cout_30_8_0;

full_adder fa_30_8_0(sum_30_8_0, cout_30_8_0, A6B24, A5B25, A4B26);

wire sum_30_9_0, cout_30_9_0;

full_adder fa_30_9_0(sum_30_9_0, cout_30_9_0, A3B27, A2B28, A1B29);

wire sum_31_0_0, cout_31_0_0;

full_adder fa_31_0_0(sum_31_0_0, cout_31_0_0, A31B0, A30B1, A29B2);

wire sum_31_1_0, cout_31_1_0;

full_adder fa_31_1_0(sum_31_1_0, cout_31_1_0, A28B3, A27B4, A26B5);

wire sum_31_2_0, cout_31_2_0;

full_adder fa_31_2_0(sum_31_2_0, cout_31_2_0, A25B6, A24B7, A23B8);

wire sum_31_3_0, cout_31_3_0;

full_adder fa_31_3_0(sum_31_3_0, cout_31_3_0, A22B9, A21B10, A20B11);

wire sum_31_4_0, cout_31_4_0;

full_adder fa_31_4_0(sum_31_4_0, cout_31_4_0, A19B12, A18B13, A17B14);

wire sum_31_5_0, cout_31_5_0;

full_adder fa_31_5_0(sum_31_5_0, cout_31_5_0, A16B15, A15B16, A14B17);

wire sum_31_6_0, cout_31_6_0;

full_adder fa_31_6_0(sum_31_6_0, cout_31_6_0, A13B18, A12B19, A11B20);

wire sum_31_7_0, cout_31_7_0;

full_adder fa_31_7_0(sum_31_7_0, cout_31_7_0, A10B21, A9B22, A8B23);

wire sum_31_8_0, cout_31_8_0;

full_adder fa_31_8_0(sum_31_8_0, cout_31_8_0, A7B24, A6B25, A5B26);

wire sum_31_9_0, cout_31_9_0;

full_adder fa_31_9_0(sum_31_9_0, cout_31_9_0, A4B27, A3B28, A2B29);

wire sum_31_10_0, cout_31_10_0;

half_adder ha_31_10_0(sum_31_10_0, cout_31_10_0, A1B30, A0B31);

wire sum_32_0_0, cout_32_0_0;

full_adder fa_32_0_0(sum_32_0_0, cout_32_0_0, A31B1, A30B2, A29B3);

wire sum_32_1_0, cout_32_1_0;

full_adder fa_32_1_0(sum_32_1_0, cout_32_1_0, A28B4, A27B5, A26B6);

wire sum_32_2_0, cout_32_2_0;

full_adder fa_32_2_0(sum_32_2_0, cout_32_2_0, A25B7, A24B8, A23B9);

wire sum_32_3_0, cout_32_3_0;

full_adder fa_32_3_0(sum_32_3_0, cout_32_3_0, A22B10, A21B11, A20B12);

wire sum_32_4_0, cout_32_4_0;

full_adder fa_32_4_0(sum_32_4_0, cout_32_4_0, A19B13, A18B14, A17B15);

wire sum_32_5_0, cout_32_5_0;

full_adder fa_32_5_0(sum_32_5_0, cout_32_5_0, A16B16, A15B17, A14B18);

wire sum_32_6_0, cout_32_6_0;

full_adder fa_32_6_0(sum_32_6_0, cout_32_6_0, A13B19, A12B20, A11B21);

wire sum_32_7_0, cout_32_7_0;

full_adder fa_32_7_0(sum_32_7_0, cout_32_7_0, A10B22, A9B23, A8B24);

wire sum_32_8_0, cout_32_8_0;

full_adder fa_32_8_0(sum_32_8_0, cout_32_8_0, A7B25, A6B26, A5B27);

wire sum_32_9_0, cout_32_9_0;

full_adder fa_32_9_0(sum_32_9_0, cout_32_9_0, A4B28, A3B29, A2B30);

wire sum_33_0_0, cout_33_0_0;

full_adder fa_33_0_0(sum_33_0_0, cout_33_0_0, A31B2, A30B3, A29B4);

wire sum_33_1_0, cout_33_1_0;

full_adder fa_33_1_0(sum_33_1_0, cout_33_1_0, A28B5, A27B6, A26B7);

wire sum_33_2_0, cout_33_2_0;

full_adder fa_33_2_0(sum_33_2_0, cout_33_2_0, A25B8, A24B9, A23B10);

wire sum_33_3_0, cout_33_3_0;

full_adder fa_33_3_0(sum_33_3_0, cout_33_3_0, A22B11, A21B12, A20B13);

wire sum_33_4_0, cout_33_4_0;

full_adder fa_33_4_0(sum_33_4_0, cout_33_4_0, A19B14, A18B15, A17B16);

wire sum_33_5_0, cout_33_5_0;

full_adder fa_33_5_0(sum_33_5_0, cout_33_5_0, A16B17, A15B18, A14B19);

wire sum_33_6_0, cout_33_6_0;

full_adder fa_33_6_0(sum_33_6_0, cout_33_6_0, A13B20, A12B21, A11B22);

wire sum_33_7_0, cout_33_7_0;

full_adder fa_33_7_0(sum_33_7_0, cout_33_7_0, A10B23, A9B24, A8B25);

wire sum_33_8_0, cout_33_8_0;

full_adder fa_33_8_0(sum_33_8_0, cout_33_8_0, A7B26, A6B27, A5B28);

wire sum_33_9_0, cout_33_9_0;

full_adder fa_33_9_0(sum_33_9_0, cout_33_9_0, A4B29, A3B30, A2B31);

wire sum_34_0_0, cout_34_0_0;

full_adder fa_34_0_0(sum_34_0_0, cout_34_0_0, A31B3, A30B4, A29B5);

wire sum_34_1_0, cout_34_1_0;

full_adder fa_34_1_0(sum_34_1_0, cout_34_1_0, A28B6, A27B7, A26B8);

wire sum_34_2_0, cout_34_2_0;

full_adder fa_34_2_0(sum_34_2_0, cout_34_2_0, A25B9, A24B10, A23B11);

wire sum_34_3_0, cout_34_3_0;

full_adder fa_34_3_0(sum_34_3_0, cout_34_3_0, A22B12, A21B13, A20B14);

wire sum_34_4_0, cout_34_4_0;

full_adder fa_34_4_0(sum_34_4_0, cout_34_4_0, A19B15, A18B16, A17B17);

wire sum_34_5_0, cout_34_5_0;

full_adder fa_34_5_0(sum_34_5_0, cout_34_5_0, A16B18, A15B19, A14B20);

wire sum_34_6_0, cout_34_6_0;

full_adder fa_34_6_0(sum_34_6_0, cout_34_6_0, A13B21, A12B22, A11B23);

wire sum_34_7_0, cout_34_7_0;

full_adder fa_34_7_0(sum_34_7_0, cout_34_7_0, A10B24, A9B25, A8B26);

wire sum_34_8_0, cout_34_8_0;

full_adder fa_34_8_0(sum_34_8_0, cout_34_8_0, A7B27, A6B28, A5B29);

wire sum_34_9_0, cout_34_9_0;

half_adder ha_34_9_0(sum_34_9_0, cout_34_9_0, A4B30, A3B31);

wire sum_35_0_0, cout_35_0_0;

full_adder fa_35_0_0(sum_35_0_0, cout_35_0_0, A31B4, A30B5, A29B6);

wire sum_35_1_0, cout_35_1_0;

full_adder fa_35_1_0(sum_35_1_0, cout_35_1_0, A28B7, A27B8, A26B9);

wire sum_35_2_0, cout_35_2_0;

full_adder fa_35_2_0(sum_35_2_0, cout_35_2_0, A25B10, A24B11, A23B12);

wire sum_35_3_0, cout_35_3_0;

full_adder fa_35_3_0(sum_35_3_0, cout_35_3_0, A22B13, A21B14, A20B15);

wire sum_35_4_0, cout_35_4_0;

full_adder fa_35_4_0(sum_35_4_0, cout_35_4_0, A19B16, A18B17, A17B18);

wire sum_35_5_0, cout_35_5_0;

full_adder fa_35_5_0(sum_35_5_0, cout_35_5_0, A16B19, A15B20, A14B21);

wire sum_35_6_0, cout_35_6_0;

full_adder fa_35_6_0(sum_35_6_0, cout_35_6_0, A13B22, A12B23, A11B24);

wire sum_35_7_0, cout_35_7_0;

full_adder fa_35_7_0(sum_35_7_0, cout_35_7_0, A10B25, A9B26, A8B27);

wire sum_35_8_0, cout_35_8_0;

full_adder fa_35_8_0(sum_35_8_0, cout_35_8_0, A7B28, A6B29, A5B30);

wire sum_36_0_0, cout_36_0_0;

full_adder fa_36_0_0(sum_36_0_0, cout_36_0_0, A31B5, A30B6, A29B7);

wire sum_36_1_0, cout_36_1_0;

full_adder fa_36_1_0(sum_36_1_0, cout_36_1_0, A28B8, A27B9, A26B10);

wire sum_36_2_0, cout_36_2_0;

full_adder fa_36_2_0(sum_36_2_0, cout_36_2_0, A25B11, A24B12, A23B13);

wire sum_36_3_0, cout_36_3_0;

full_adder fa_36_3_0(sum_36_3_0, cout_36_3_0, A22B14, A21B15, A20B16);

wire sum_36_4_0, cout_36_4_0;

full_adder fa_36_4_0(sum_36_4_0, cout_36_4_0, A19B17, A18B18, A17B19);

wire sum_36_5_0, cout_36_5_0;

full_adder fa_36_5_0(sum_36_5_0, cout_36_5_0, A16B20, A15B21, A14B22);

wire sum_36_6_0, cout_36_6_0;

full_adder fa_36_6_0(sum_36_6_0, cout_36_6_0, A13B23, A12B24, A11B25);

wire sum_36_7_0, cout_36_7_0;

full_adder fa_36_7_0(sum_36_7_0, cout_36_7_0, A10B26, A9B27, A8B28);

wire sum_36_8_0, cout_36_8_0;

full_adder fa_36_8_0(sum_36_8_0, cout_36_8_0, A7B29, A6B30, A5B31);

wire sum_37_0_0, cout_37_0_0;

full_adder fa_37_0_0(sum_37_0_0, cout_37_0_0, A31B6, A30B7, A29B8);

wire sum_37_1_0, cout_37_1_0;

full_adder fa_37_1_0(sum_37_1_0, cout_37_1_0, A28B9, A27B10, A26B11);

wire sum_37_2_0, cout_37_2_0;

full_adder fa_37_2_0(sum_37_2_0, cout_37_2_0, A25B12, A24B13, A23B14);

wire sum_37_3_0, cout_37_3_0;

full_adder fa_37_3_0(sum_37_3_0, cout_37_3_0, A22B15, A21B16, A20B17);

wire sum_37_4_0, cout_37_4_0;

full_adder fa_37_4_0(sum_37_4_0, cout_37_4_0, A19B18, A18B19, A17B20);

wire sum_37_5_0, cout_37_5_0;

full_adder fa_37_5_0(sum_37_5_0, cout_37_5_0, A16B21, A15B22, A14B23);

wire sum_37_6_0, cout_37_6_0;

full_adder fa_37_6_0(sum_37_6_0, cout_37_6_0, A13B24, A12B25, A11B26);

wire sum_37_7_0, cout_37_7_0;

full_adder fa_37_7_0(sum_37_7_0, cout_37_7_0, A10B27, A9B28, A8B29);

wire sum_37_8_0, cout_37_8_0;

half_adder ha_37_8_0(sum_37_8_0, cout_37_8_0, A7B30, A6B31);

wire sum_38_0_0, cout_38_0_0;

full_adder fa_38_0_0(sum_38_0_0, cout_38_0_0, A31B7, A30B8, A29B9);

wire sum_38_1_0, cout_38_1_0;

full_adder fa_38_1_0(sum_38_1_0, cout_38_1_0, A28B10, A27B11, A26B12);

wire sum_38_2_0, cout_38_2_0;

full_adder fa_38_2_0(sum_38_2_0, cout_38_2_0, A25B13, A24B14, A23B15);

wire sum_38_3_0, cout_38_3_0;

full_adder fa_38_3_0(sum_38_3_0, cout_38_3_0, A22B16, A21B17, A20B18);

wire sum_38_4_0, cout_38_4_0;

full_adder fa_38_4_0(sum_38_4_0, cout_38_4_0, A19B19, A18B20, A17B21);

wire sum_38_5_0, cout_38_5_0;

full_adder fa_38_5_0(sum_38_5_0, cout_38_5_0, A16B22, A15B23, A14B24);

wire sum_38_6_0, cout_38_6_0;

full_adder fa_38_6_0(sum_38_6_0, cout_38_6_0, A13B25, A12B26, A11B27);

wire sum_38_7_0, cout_38_7_0;

full_adder fa_38_7_0(sum_38_7_0, cout_38_7_0, A10B28, A9B29, A8B30);

wire sum_39_0_0, cout_39_0_0;

full_adder fa_39_0_0(sum_39_0_0, cout_39_0_0, A31B8, A30B9, A29B10);

wire sum_39_1_0, cout_39_1_0;

full_adder fa_39_1_0(sum_39_1_0, cout_39_1_0, A28B11, A27B12, A26B13);

wire sum_39_2_0, cout_39_2_0;

full_adder fa_39_2_0(sum_39_2_0, cout_39_2_0, A25B14, A24B15, A23B16);

wire sum_39_3_0, cout_39_3_0;

full_adder fa_39_3_0(sum_39_3_0, cout_39_3_0, A22B17, A21B18, A20B19);

wire sum_39_4_0, cout_39_4_0;

full_adder fa_39_4_0(sum_39_4_0, cout_39_4_0, A19B20, A18B21, A17B22);

wire sum_39_5_0, cout_39_5_0;

full_adder fa_39_5_0(sum_39_5_0, cout_39_5_0, A16B23, A15B24, A14B25);

wire sum_39_6_0, cout_39_6_0;

full_adder fa_39_6_0(sum_39_6_0, cout_39_6_0, A13B26, A12B27, A11B28);

wire sum_39_7_0, cout_39_7_0;

full_adder fa_39_7_0(sum_39_7_0, cout_39_7_0, A10B29, A9B30, A8B31);

wire sum_40_0_0, cout_40_0_0;

full_adder fa_40_0_0(sum_40_0_0, cout_40_0_0, A31B9, A30B10, A29B11);

wire sum_40_1_0, cout_40_1_0;

full_adder fa_40_1_0(sum_40_1_0, cout_40_1_0, A28B12, A27B13, A26B14);

wire sum_40_2_0, cout_40_2_0;

full_adder fa_40_2_0(sum_40_2_0, cout_40_2_0, A25B15, A24B16, A23B17);

wire sum_40_3_0, cout_40_3_0;

full_adder fa_40_3_0(sum_40_3_0, cout_40_3_0, A22B18, A21B19, A20B20);

wire sum_40_4_0, cout_40_4_0;

full_adder fa_40_4_0(sum_40_4_0, cout_40_4_0, A19B21, A18B22, A17B23);

wire sum_40_5_0, cout_40_5_0;

full_adder fa_40_5_0(sum_40_5_0, cout_40_5_0, A16B24, A15B25, A14B26);

wire sum_40_6_0, cout_40_6_0;

full_adder fa_40_6_0(sum_40_6_0, cout_40_6_0, A13B27, A12B28, A11B29);

wire sum_40_7_0, cout_40_7_0;

half_adder ha_40_7_0(sum_40_7_0, cout_40_7_0, A10B30, A9B31);

wire sum_41_0_0, cout_41_0_0;

full_adder fa_41_0_0(sum_41_0_0, cout_41_0_0, A31B10, A30B11, A29B12);

wire sum_41_1_0, cout_41_1_0;

full_adder fa_41_1_0(sum_41_1_0, cout_41_1_0, A28B13, A27B14, A26B15);

wire sum_41_2_0, cout_41_2_0;

full_adder fa_41_2_0(sum_41_2_0, cout_41_2_0, A25B16, A24B17, A23B18);

wire sum_41_3_0, cout_41_3_0;

full_adder fa_41_3_0(sum_41_3_0, cout_41_3_0, A22B19, A21B20, A20B21);

wire sum_41_4_0, cout_41_4_0;

full_adder fa_41_4_0(sum_41_4_0, cout_41_4_0, A19B22, A18B23, A17B24);

wire sum_41_5_0, cout_41_5_0;

full_adder fa_41_5_0(sum_41_5_0, cout_41_5_0, A16B25, A15B26, A14B27);

wire sum_41_6_0, cout_41_6_0;

full_adder fa_41_6_0(sum_41_6_0, cout_41_6_0, A13B28, A12B29, A11B30);

wire sum_42_0_0, cout_42_0_0;

full_adder fa_42_0_0(sum_42_0_0, cout_42_0_0, A31B11, A30B12, A29B13);

wire sum_42_1_0, cout_42_1_0;

full_adder fa_42_1_0(sum_42_1_0, cout_42_1_0, A28B14, A27B15, A26B16);

wire sum_42_2_0, cout_42_2_0;

full_adder fa_42_2_0(sum_42_2_0, cout_42_2_0, A25B17, A24B18, A23B19);

wire sum_42_3_0, cout_42_3_0;

full_adder fa_42_3_0(sum_42_3_0, cout_42_3_0, A22B20, A21B21, A20B22);

wire sum_42_4_0, cout_42_4_0;

full_adder fa_42_4_0(sum_42_4_0, cout_42_4_0, A19B23, A18B24, A17B25);

wire sum_42_5_0, cout_42_5_0;

full_adder fa_42_5_0(sum_42_5_0, cout_42_5_0, A16B26, A15B27, A14B28);

wire sum_42_6_0, cout_42_6_0;

full_adder fa_42_6_0(sum_42_6_0, cout_42_6_0, A13B29, A12B30, A11B31);

wire sum_43_0_0, cout_43_0_0;

full_adder fa_43_0_0(sum_43_0_0, cout_43_0_0, A31B12, A30B13, A29B14);

wire sum_43_1_0, cout_43_1_0;

full_adder fa_43_1_0(sum_43_1_0, cout_43_1_0, A28B15, A27B16, A26B17);

wire sum_43_2_0, cout_43_2_0;

full_adder fa_43_2_0(sum_43_2_0, cout_43_2_0, A25B18, A24B19, A23B20);

wire sum_43_3_0, cout_43_3_0;

full_adder fa_43_3_0(sum_43_3_0, cout_43_3_0, A22B21, A21B22, A20B23);

wire sum_43_4_0, cout_43_4_0;

full_adder fa_43_4_0(sum_43_4_0, cout_43_4_0, A19B24, A18B25, A17B26);

wire sum_43_5_0, cout_43_5_0;

full_adder fa_43_5_0(sum_43_5_0, cout_43_5_0, A16B27, A15B28, A14B29);

wire sum_43_6_0, cout_43_6_0;

half_adder ha_43_6_0(sum_43_6_0, cout_43_6_0, A13B30, A12B31);

wire sum_44_0_0, cout_44_0_0;

full_adder fa_44_0_0(sum_44_0_0, cout_44_0_0, A31B13, A30B14, A29B15);

wire sum_44_1_0, cout_44_1_0;

full_adder fa_44_1_0(sum_44_1_0, cout_44_1_0, A28B16, A27B17, A26B18);

wire sum_44_2_0, cout_44_2_0;

full_adder fa_44_2_0(sum_44_2_0, cout_44_2_0, A25B19, A24B20, A23B21);

wire sum_44_3_0, cout_44_3_0;

full_adder fa_44_3_0(sum_44_3_0, cout_44_3_0, A22B22, A21B23, A20B24);

wire sum_44_4_0, cout_44_4_0;

full_adder fa_44_4_0(sum_44_4_0, cout_44_4_0, A19B25, A18B26, A17B27);

wire sum_44_5_0, cout_44_5_0;

full_adder fa_44_5_0(sum_44_5_0, cout_44_5_0, A16B28, A15B29, A14B30);

wire sum_45_0_0, cout_45_0_0;

full_adder fa_45_0_0(sum_45_0_0, cout_45_0_0, A31B14, A30B15, A29B16);

wire sum_45_1_0, cout_45_1_0;

full_adder fa_45_1_0(sum_45_1_0, cout_45_1_0, A28B17, A27B18, A26B19);

wire sum_45_2_0, cout_45_2_0;

full_adder fa_45_2_0(sum_45_2_0, cout_45_2_0, A25B20, A24B21, A23B22);

wire sum_45_3_0, cout_45_3_0;

full_adder fa_45_3_0(sum_45_3_0, cout_45_3_0, A22B23, A21B24, A20B25);

wire sum_45_4_0, cout_45_4_0;

full_adder fa_45_4_0(sum_45_4_0, cout_45_4_0, A19B26, A18B27, A17B28);

wire sum_45_5_0, cout_45_5_0;

full_adder fa_45_5_0(sum_45_5_0, cout_45_5_0, A16B29, A15B30, A14B31);

wire sum_46_0_0, cout_46_0_0;

full_adder fa_46_0_0(sum_46_0_0, cout_46_0_0, A31B15, A30B16, A29B17);

wire sum_46_1_0, cout_46_1_0;

full_adder fa_46_1_0(sum_46_1_0, cout_46_1_0, A28B18, A27B19, A26B20);

wire sum_46_2_0, cout_46_2_0;

full_adder fa_46_2_0(sum_46_2_0, cout_46_2_0, A25B21, A24B22, A23B23);

wire sum_46_3_0, cout_46_3_0;

full_adder fa_46_3_0(sum_46_3_0, cout_46_3_0, A22B24, A21B25, A20B26);

wire sum_46_4_0, cout_46_4_0;

full_adder fa_46_4_0(sum_46_4_0, cout_46_4_0, A19B27, A18B28, A17B29);

wire sum_46_5_0, cout_46_5_0;

half_adder ha_46_5_0(sum_46_5_0, cout_46_5_0, A16B30, A15B31);

wire sum_47_0_0, cout_47_0_0;

full_adder fa_47_0_0(sum_47_0_0, cout_47_0_0, A31B16, A30B17, A29B18);

wire sum_47_1_0, cout_47_1_0;

full_adder fa_47_1_0(sum_47_1_0, cout_47_1_0, A28B19, A27B20, A26B21);

wire sum_47_2_0, cout_47_2_0;

full_adder fa_47_2_0(sum_47_2_0, cout_47_2_0, A25B22, A24B23, A23B24);

wire sum_47_3_0, cout_47_3_0;

full_adder fa_47_3_0(sum_47_3_0, cout_47_3_0, A22B25, A21B26, A20B27);

wire sum_47_4_0, cout_47_4_0;

full_adder fa_47_4_0(sum_47_4_0, cout_47_4_0, A19B28, A18B29, A17B30);

wire sum_48_0_0, cout_48_0_0;

full_adder fa_48_0_0(sum_48_0_0, cout_48_0_0, A31B17, A30B18, A29B19);

wire sum_48_1_0, cout_48_1_0;

full_adder fa_48_1_0(sum_48_1_0, cout_48_1_0, A28B20, A27B21, A26B22);

wire sum_48_2_0, cout_48_2_0;

full_adder fa_48_2_0(sum_48_2_0, cout_48_2_0, A25B23, A24B24, A23B25);

wire sum_48_3_0, cout_48_3_0;

full_adder fa_48_3_0(sum_48_3_0, cout_48_3_0, A22B26, A21B27, A20B28);

wire sum_48_4_0, cout_48_4_0;

full_adder fa_48_4_0(sum_48_4_0, cout_48_4_0, A19B29, A18B30, A17B31);

wire sum_49_0_0, cout_49_0_0;

full_adder fa_49_0_0(sum_49_0_0, cout_49_0_0, A31B18, A30B19, A29B20);

wire sum_49_1_0, cout_49_1_0;

full_adder fa_49_1_0(sum_49_1_0, cout_49_1_0, A28B21, A27B22, A26B23);

wire sum_49_2_0, cout_49_2_0;

full_adder fa_49_2_0(sum_49_2_0, cout_49_2_0, A25B24, A24B25, A23B26);

wire sum_49_3_0, cout_49_3_0;

full_adder fa_49_3_0(sum_49_3_0, cout_49_3_0, A22B27, A21B28, A20B29);

wire sum_49_4_0, cout_49_4_0;

half_adder ha_49_4_0(sum_49_4_0, cout_49_4_0, A19B30, A18B31);

wire sum_50_0_0, cout_50_0_0;

full_adder fa_50_0_0(sum_50_0_0, cout_50_0_0, A31B19, A30B20, A29B21);

wire sum_50_1_0, cout_50_1_0;

full_adder fa_50_1_0(sum_50_1_0, cout_50_1_0, A28B22, A27B23, A26B24);

wire sum_50_2_0, cout_50_2_0;

full_adder fa_50_2_0(sum_50_2_0, cout_50_2_0, A25B25, A24B26, A23B27);

wire sum_50_3_0, cout_50_3_0;

full_adder fa_50_3_0(sum_50_3_0, cout_50_3_0, A22B28, A21B29, A20B30);

wire sum_51_0_0, cout_51_0_0;

full_adder fa_51_0_0(sum_51_0_0, cout_51_0_0, A31B20, A30B21, A29B22);

wire sum_51_1_0, cout_51_1_0;

full_adder fa_51_1_0(sum_51_1_0, cout_51_1_0, A28B23, A27B24, A26B25);

wire sum_51_2_0, cout_51_2_0;

full_adder fa_51_2_0(sum_51_2_0, cout_51_2_0, A25B26, A24B27, A23B28);

wire sum_51_3_0, cout_51_3_0;

full_adder fa_51_3_0(sum_51_3_0, cout_51_3_0, A22B29, A21B30, A20B31);

wire sum_52_0_0, cout_52_0_0;

full_adder fa_52_0_0(sum_52_0_0, cout_52_0_0, A31B21, A30B22, A29B23);

wire sum_52_1_0, cout_52_1_0;

full_adder fa_52_1_0(sum_52_1_0, cout_52_1_0, A28B24, A27B25, A26B26);

wire sum_52_2_0, cout_52_2_0;

full_adder fa_52_2_0(sum_52_2_0, cout_52_2_0, A25B27, A24B28, A23B29);

wire sum_52_3_0, cout_52_3_0;

half_adder ha_52_3_0(sum_52_3_0, cout_52_3_0, A22B30, A21B31);

wire sum_53_0_0, cout_53_0_0;

full_adder fa_53_0_0(sum_53_0_0, cout_53_0_0, A31B22, A30B23, A29B24);

wire sum_53_1_0, cout_53_1_0;

full_adder fa_53_1_0(sum_53_1_0, cout_53_1_0, A28B25, A27B26, A26B27);

wire sum_53_2_0, cout_53_2_0;

full_adder fa_53_2_0(sum_53_2_0, cout_53_2_0, A25B28, A24B29, A23B30);

wire sum_54_0_0, cout_54_0_0;

full_adder fa_54_0_0(sum_54_0_0, cout_54_0_0, A31B23, A30B24, A29B25);

wire sum_54_1_0, cout_54_1_0;

full_adder fa_54_1_0(sum_54_1_0, cout_54_1_0, A28B26, A27B27, A26B28);

wire sum_54_2_0, cout_54_2_0;

full_adder fa_54_2_0(sum_54_2_0, cout_54_2_0, A25B29, A24B30, A23B31);

wire sum_55_0_0, cout_55_0_0;

full_adder fa_55_0_0(sum_55_0_0, cout_55_0_0, A31B24, A30B25, A29B26);

wire sum_55_1_0, cout_55_1_0;

full_adder fa_55_1_0(sum_55_1_0, cout_55_1_0, A28B27, A27B28, A26B29);

wire sum_55_2_0, cout_55_2_0;

half_adder ha_55_2_0(sum_55_2_0, cout_55_2_0, A25B30, A24B31);

wire sum_56_0_0, cout_56_0_0;

full_adder fa_56_0_0(sum_56_0_0, cout_56_0_0, A31B25, A30B26, A29B27);

wire sum_56_1_0, cout_56_1_0;

full_adder fa_56_1_0(sum_56_1_0, cout_56_1_0, A28B28, A27B29, A26B30);

wire sum_57_0_0, cout_57_0_0;

full_adder fa_57_0_0(sum_57_0_0, cout_57_0_0, A31B26, A30B27, A29B28);

wire sum_57_1_0, cout_57_1_0;

full_adder fa_57_1_0(sum_57_1_0, cout_57_1_0, A28B29, A27B30, A26B31);

wire sum_58_0_0, cout_58_0_0;

full_adder fa_58_0_0(sum_58_0_0, cout_58_0_0, A31B27, A30B28, A29B29);

wire sum_58_1_0, cout_58_1_0;

half_adder ha_58_1_0(sum_58_1_0, cout_58_1_0, A28B30, A27B31);

wire sum_59_0_0, cout_59_0_0;

full_adder fa_59_0_0(sum_59_0_0, cout_59_0_0, A31B28, A30B29, A29B30);

wire sum_60_0_0, cout_60_0_0;

full_adder fa_60_0_0(sum_60_0_0, cout_60_0_0, A31B29, A30B30, A29B31);

wire sum_3_0_1, cout_3_0_1;

half_adder ha_3_0_1(sum_3_0_1, cout_3_0_1, A0B3, cout_2_0_0);

wire sum_4_0_1, cout_4_0_1;

full_adder fa_4_0_1(sum_4_0_1, cout_4_0_1, cout_3_0_0, sum_4_0_0, sum_4_1_0);

wire sum_5_0_1, cout_5_0_1;

full_adder fa_5_0_1(sum_5_0_1, cout_5_0_1, cout_4_0_0, cout_4_1_0, sum_5_0_0);

wire sum_6_0_1, cout_6_0_1;

full_adder fa_6_0_1(sum_6_0_1, cout_6_0_1, A0B6, cout_5_0_0, cout_5_1_0);

wire sum_6_1_1, cout_6_1_1;

half_adder ha_6_1_1(sum_6_1_1, cout_6_1_1, sum_6_0_0, sum_6_1_0);

wire sum_7_0_1, cout_7_0_1;

full_adder fa_7_0_1(sum_7_0_1, cout_7_0_1, cout_6_0_0, cout_6_1_0, sum_7_0_0);

wire sum_7_1_1, cout_7_1_1;

half_adder ha_7_1_1(sum_7_1_1, cout_7_1_1, sum_7_1_0, sum_7_2_0);

wire sum_8_0_1, cout_8_0_1;

full_adder fa_8_0_1(sum_8_0_1, cout_8_0_1, cout_7_0_0, cout_7_1_0, cout_7_2_0);

wire sum_8_1_1, cout_8_1_1;

full_adder fa_8_1_1(sum_8_1_1, cout_8_1_1, sum_8_0_0, sum_8_1_0, sum_8_2_0);

wire sum_9_0_1, cout_9_0_1;

full_adder fa_9_0_1(sum_9_0_1, cout_9_0_1, A0B9, cout_8_0_0, cout_8_1_0);

wire sum_9_1_1, cout_9_1_1;

full_adder fa_9_1_1(sum_9_1_1, cout_9_1_1, cout_8_2_0, sum_9_0_0, sum_9_1_0);

wire sum_10_0_1, cout_10_0_1;

full_adder fa_10_0_1(sum_10_0_1, cout_10_0_1, cout_9_0_0, cout_9_1_0, cout_9_2_0);

wire sum_10_1_1, cout_10_1_1;

full_adder fa_10_1_1(sum_10_1_1, cout_10_1_1, sum_10_0_0, sum_10_1_0, sum_10_2_0);

wire sum_11_0_1, cout_11_0_1;

full_adder fa_11_0_1(sum_11_0_1, cout_11_0_1, cout_10_0_0, cout_10_1_0, cout_10_2_0);

wire sum_11_1_1, cout_11_1_1;

full_adder fa_11_1_1(sum_11_1_1, cout_11_1_1, cout_10_3_0, sum_11_0_0, sum_11_1_0);

wire sum_11_2_1, cout_11_2_1;

half_adder ha_11_2_1(sum_11_2_1, cout_11_2_1, sum_11_2_0, sum_11_3_0);

wire sum_12_0_1, cout_12_0_1;

full_adder fa_12_0_1(sum_12_0_1, cout_12_0_1, A0B12, cout_11_0_0, cout_11_1_0);

wire sum_12_1_1, cout_12_1_1;

full_adder fa_12_1_1(sum_12_1_1, cout_12_1_1, cout_11_2_0, cout_11_3_0, sum_12_0_0);

wire sum_12_2_1, cout_12_2_1;

full_adder fa_12_2_1(sum_12_2_1, cout_12_2_1, sum_12_1_0, sum_12_2_0, sum_12_3_0);

wire sum_13_0_1, cout_13_0_1;

full_adder fa_13_0_1(sum_13_0_1, cout_13_0_1, cout_12_0_0, cout_12_1_0, cout_12_2_0);

wire sum_13_1_1, cout_13_1_1;

full_adder fa_13_1_1(sum_13_1_1, cout_13_1_1, cout_12_3_0, sum_13_0_0, sum_13_1_0);

wire sum_13_2_1, cout_13_2_1;

full_adder fa_13_2_1(sum_13_2_1, cout_13_2_1, sum_13_2_0, sum_13_3_0, sum_13_4_0);

wire sum_14_0_1, cout_14_0_1;

full_adder fa_14_0_1(sum_14_0_1, cout_14_0_1, cout_13_0_0, cout_13_1_0, cout_13_2_0);

wire sum_14_1_1, cout_14_1_1;

full_adder fa_14_1_1(sum_14_1_1, cout_14_1_1, cout_13_3_0, cout_13_4_0, sum_14_0_0);

wire sum_14_2_1, cout_14_2_1;

full_adder fa_14_2_1(sum_14_2_1, cout_14_2_1, sum_14_1_0, sum_14_2_0, sum_14_3_0);

wire sum_15_0_1, cout_15_0_1;

full_adder fa_15_0_1(sum_15_0_1, cout_15_0_1, A0B15, cout_14_0_0, cout_14_1_0);

wire sum_15_1_1, cout_15_1_1;

full_adder fa_15_1_1(sum_15_1_1, cout_15_1_1, cout_14_2_0, cout_14_3_0, cout_14_4_0);

wire sum_15_2_1, cout_15_2_1;

full_adder fa_15_2_1(sum_15_2_1, cout_15_2_1, sum_15_0_0, sum_15_1_0, sum_15_2_0);

wire sum_15_3_1, cout_15_3_1;

half_adder ha_15_3_1(sum_15_3_1, cout_15_3_1, sum_15_3_0, sum_15_4_0);

wire sum_16_0_1, cout_16_0_1;

full_adder fa_16_0_1(sum_16_0_1, cout_16_0_1, cout_15_0_0, cout_15_1_0, cout_15_2_0);

wire sum_16_1_1, cout_16_1_1;

full_adder fa_16_1_1(sum_16_1_1, cout_16_1_1, cout_15_3_0, cout_15_4_0, sum_16_0_0);

wire sum_16_2_1, cout_16_2_1;

full_adder fa_16_2_1(sum_16_2_1, cout_16_2_1, sum_16_1_0, sum_16_2_0, sum_16_3_0);

wire sum_16_3_1, cout_16_3_1;

half_adder ha_16_3_1(sum_16_3_1, cout_16_3_1, sum_16_4_0, sum_16_5_0);

wire sum_17_0_1, cout_17_0_1;

full_adder fa_17_0_1(sum_17_0_1, cout_17_0_1, cout_16_0_0, cout_16_1_0, cout_16_2_0);

wire sum_17_1_1, cout_17_1_1;

full_adder fa_17_1_1(sum_17_1_1, cout_17_1_1, cout_16_3_0, cout_16_4_0, cout_16_5_0);

wire sum_17_2_1, cout_17_2_1;

full_adder fa_17_2_1(sum_17_2_1, cout_17_2_1, sum_17_0_0, sum_17_1_0, sum_17_2_0);

wire sum_17_3_1, cout_17_3_1;

full_adder fa_17_3_1(sum_17_3_1, cout_17_3_1, sum_17_3_0, sum_17_4_0, sum_17_5_0);

wire sum_18_0_1, cout_18_0_1;

full_adder fa_18_0_1(sum_18_0_1, cout_18_0_1, A0B18, cout_17_0_0, cout_17_1_0);

wire sum_18_1_1, cout_18_1_1;

full_adder fa_18_1_1(sum_18_1_1, cout_18_1_1, cout_17_2_0, cout_17_3_0, cout_17_4_0);

wire sum_18_2_1, cout_18_2_1;

full_adder fa_18_2_1(sum_18_2_1, cout_18_2_1, cout_17_5_0, sum_18_0_0, sum_18_1_0);

wire sum_18_3_1, cout_18_3_1;

full_adder fa_18_3_1(sum_18_3_1, cout_18_3_1, sum_18_2_0, sum_18_3_0, sum_18_4_0);

wire sum_19_0_1, cout_19_0_1;

full_adder fa_19_0_1(sum_19_0_1, cout_19_0_1, cout_18_0_0, cout_18_1_0, cout_18_2_0);

wire sum_19_1_1, cout_19_1_1;

full_adder fa_19_1_1(sum_19_1_1, cout_19_1_1, cout_18_3_0, cout_18_4_0, cout_18_5_0);

wire sum_19_2_1, cout_19_2_1;

full_adder fa_19_2_1(sum_19_2_1, cout_19_2_1, sum_19_0_0, sum_19_1_0, sum_19_2_0);

wire sum_19_3_1, cout_19_3_1;

full_adder fa_19_3_1(sum_19_3_1, cout_19_3_1, sum_19_3_0, sum_19_4_0, sum_19_5_0);

wire sum_20_0_1, cout_20_0_1;

full_adder fa_20_0_1(sum_20_0_1, cout_20_0_1, cout_19_0_0, cout_19_1_0, cout_19_2_0);

wire sum_20_1_1, cout_20_1_1;

full_adder fa_20_1_1(sum_20_1_1, cout_20_1_1, cout_19_3_0, cout_19_4_0, cout_19_5_0);

wire sum_20_2_1, cout_20_2_1;

full_adder fa_20_2_1(sum_20_2_1, cout_20_2_1, cout_19_6_0, sum_20_0_0, sum_20_1_0);

wire sum_20_3_1, cout_20_3_1;

full_adder fa_20_3_1(sum_20_3_1, cout_20_3_1, sum_20_2_0, sum_20_3_0, sum_20_4_0);

wire sum_20_4_1, cout_20_4_1;

half_adder ha_20_4_1(sum_20_4_1, cout_20_4_1, sum_20_5_0, sum_20_6_0);

wire sum_21_0_1, cout_21_0_1;

full_adder fa_21_0_1(sum_21_0_1, cout_21_0_1, A0B21, cout_20_0_0, cout_20_1_0);

wire sum_21_1_1, cout_21_1_1;

full_adder fa_21_1_1(sum_21_1_1, cout_21_1_1, cout_20_2_0, cout_20_3_0, cout_20_4_0);

wire sum_21_2_1, cout_21_2_1;

full_adder fa_21_2_1(sum_21_2_1, cout_21_2_1, cout_20_5_0, cout_20_6_0, sum_21_0_0);

wire sum_21_3_1, cout_21_3_1;

full_adder fa_21_3_1(sum_21_3_1, cout_21_3_1, sum_21_1_0, sum_21_2_0, sum_21_3_0);

wire sum_21_4_1, cout_21_4_1;

full_adder fa_21_4_1(sum_21_4_1, cout_21_4_1, sum_21_4_0, sum_21_5_0, sum_21_6_0);

wire sum_22_0_1, cout_22_0_1;

full_adder fa_22_0_1(sum_22_0_1, cout_22_0_1, cout_21_0_0, cout_21_1_0, cout_21_2_0);

wire sum_22_1_1, cout_22_1_1;

full_adder fa_22_1_1(sum_22_1_1, cout_22_1_1, cout_21_3_0, cout_21_4_0, cout_21_5_0);

wire sum_22_2_1, cout_22_2_1;

full_adder fa_22_2_1(sum_22_2_1, cout_22_2_1, cout_21_6_0, sum_22_0_0, sum_22_1_0);

wire sum_22_3_1, cout_22_3_1;

full_adder fa_22_3_1(sum_22_3_1, cout_22_3_1, sum_22_2_0, sum_22_3_0, sum_22_4_0);

wire sum_22_4_1, cout_22_4_1;

full_adder fa_22_4_1(sum_22_4_1, cout_22_4_1, sum_22_5_0, sum_22_6_0, sum_22_7_0);

wire sum_23_0_1, cout_23_0_1;

full_adder fa_23_0_1(sum_23_0_1, cout_23_0_1, cout_22_0_0, cout_22_1_0, cout_22_2_0);

wire sum_23_1_1, cout_23_1_1;

full_adder fa_23_1_1(sum_23_1_1, cout_23_1_1, cout_22_3_0, cout_22_4_0, cout_22_5_0);

wire sum_23_2_1, cout_23_2_1;

full_adder fa_23_2_1(sum_23_2_1, cout_23_2_1, cout_22_6_0, cout_22_7_0, sum_23_0_0);

wire sum_23_3_1, cout_23_3_1;

full_adder fa_23_3_1(sum_23_3_1, cout_23_3_1, sum_23_1_0, sum_23_2_0, sum_23_3_0);

wire sum_23_4_1, cout_23_4_1;

full_adder fa_23_4_1(sum_23_4_1, cout_23_4_1, sum_23_4_0, sum_23_5_0, sum_23_6_0);

wire sum_24_0_1, cout_24_0_1;

full_adder fa_24_0_1(sum_24_0_1, cout_24_0_1, A0B24, cout_23_0_0, cout_23_1_0);

wire sum_24_1_1, cout_24_1_1;

full_adder fa_24_1_1(sum_24_1_1, cout_24_1_1, cout_23_2_0, cout_23_3_0, cout_23_4_0);

wire sum_24_2_1, cout_24_2_1;

full_adder fa_24_2_1(sum_24_2_1, cout_24_2_1, cout_23_5_0, cout_23_6_0, cout_23_7_0);

wire sum_24_3_1, cout_24_3_1;

full_adder fa_24_3_1(sum_24_3_1, cout_24_3_1, sum_24_0_0, sum_24_1_0, sum_24_2_0);

wire sum_24_4_1, cout_24_4_1;

full_adder fa_24_4_1(sum_24_4_1, cout_24_4_1, sum_24_3_0, sum_24_4_0, sum_24_5_0);

wire sum_24_5_1, cout_24_5_1;

half_adder ha_24_5_1(sum_24_5_1, cout_24_5_1, sum_24_6_0, sum_24_7_0);

wire sum_25_0_1, cout_25_0_1;

full_adder fa_25_0_1(sum_25_0_1, cout_25_0_1, cout_24_0_0, cout_24_1_0, cout_24_2_0);

wire sum_25_1_1, cout_25_1_1;

full_adder fa_25_1_1(sum_25_1_1, cout_25_1_1, cout_24_3_0, cout_24_4_0, cout_24_5_0);

wire sum_25_2_1, cout_25_2_1;

full_adder fa_25_2_1(sum_25_2_1, cout_25_2_1, cout_24_6_0, cout_24_7_0, sum_25_0_0);

wire sum_25_3_1, cout_25_3_1;

full_adder fa_25_3_1(sum_25_3_1, cout_25_3_1, sum_25_1_0, sum_25_2_0, sum_25_3_0);

wire sum_25_4_1, cout_25_4_1;

full_adder fa_25_4_1(sum_25_4_1, cout_25_4_1, sum_25_4_0, sum_25_5_0, sum_25_6_0);

wire sum_25_5_1, cout_25_5_1;

half_adder ha_25_5_1(sum_25_5_1, cout_25_5_1, sum_25_7_0, sum_25_8_0);

wire sum_26_0_1, cout_26_0_1;

full_adder fa_26_0_1(sum_26_0_1, cout_26_0_1, cout_25_0_0, cout_25_1_0, cout_25_2_0);

wire sum_26_1_1, cout_26_1_1;

full_adder fa_26_1_1(sum_26_1_1, cout_26_1_1, cout_25_3_0, cout_25_4_0, cout_25_5_0);

wire sum_26_2_1, cout_26_2_1;

full_adder fa_26_2_1(sum_26_2_1, cout_26_2_1, cout_25_6_0, cout_25_7_0, cout_25_8_0);

wire sum_26_3_1, cout_26_3_1;

full_adder fa_26_3_1(sum_26_3_1, cout_26_3_1, sum_26_0_0, sum_26_1_0, sum_26_2_0);

wire sum_26_4_1, cout_26_4_1;

full_adder fa_26_4_1(sum_26_4_1, cout_26_4_1, sum_26_3_0, sum_26_4_0, sum_26_5_0);

wire sum_26_5_1, cout_26_5_1;

full_adder fa_26_5_1(sum_26_5_1, cout_26_5_1, sum_26_6_0, sum_26_7_0, sum_26_8_0);

wire sum_27_0_1, cout_27_0_1;

full_adder fa_27_0_1(sum_27_0_1, cout_27_0_1, A0B27, cout_26_0_0, cout_26_1_0);

wire sum_27_1_1, cout_27_1_1;

full_adder fa_27_1_1(sum_27_1_1, cout_27_1_1, cout_26_2_0, cout_26_3_0, cout_26_4_0);

wire sum_27_2_1, cout_27_2_1;

full_adder fa_27_2_1(sum_27_2_1, cout_27_2_1, cout_26_5_0, cout_26_6_0, cout_26_7_0);

wire sum_27_3_1, cout_27_3_1;

full_adder fa_27_3_1(sum_27_3_1, cout_27_3_1, cout_26_8_0, sum_27_0_0, sum_27_1_0);

wire sum_27_4_1, cout_27_4_1;

full_adder fa_27_4_1(sum_27_4_1, cout_27_4_1, sum_27_2_0, sum_27_3_0, sum_27_4_0);

wire sum_27_5_1, cout_27_5_1;

full_adder fa_27_5_1(sum_27_5_1, cout_27_5_1, sum_27_5_0, sum_27_6_0, sum_27_7_0);

wire sum_28_0_1, cout_28_0_1;

full_adder fa_28_0_1(sum_28_0_1, cout_28_0_1, cout_27_0_0, cout_27_1_0, cout_27_2_0);

wire sum_28_1_1, cout_28_1_1;

full_adder fa_28_1_1(sum_28_1_1, cout_28_1_1, cout_27_3_0, cout_27_4_0, cout_27_5_0);

wire sum_28_2_1, cout_28_2_1;

full_adder fa_28_2_1(sum_28_2_1, cout_28_2_1, cout_27_6_0, cout_27_7_0, cout_27_8_0);

wire sum_28_3_1, cout_28_3_1;

full_adder fa_28_3_1(sum_28_3_1, cout_28_3_1, sum_28_0_0, sum_28_1_0, sum_28_2_0);

wire sum_28_4_1, cout_28_4_1;

full_adder fa_28_4_1(sum_28_4_1, cout_28_4_1, sum_28_3_0, sum_28_4_0, sum_28_5_0);

wire sum_28_5_1, cout_28_5_1;

full_adder fa_28_5_1(sum_28_5_1, cout_28_5_1, sum_28_6_0, sum_28_7_0, sum_28_8_0);

wire sum_29_0_1, cout_29_0_1;

full_adder fa_29_0_1(sum_29_0_1, cout_29_0_1, cout_28_0_0, cout_28_1_0, cout_28_2_0);

wire sum_29_1_1, cout_29_1_1;

full_adder fa_29_1_1(sum_29_1_1, cout_29_1_1, cout_28_3_0, cout_28_4_0, cout_28_5_0);

wire sum_29_2_1, cout_29_2_1;

full_adder fa_29_2_1(sum_29_2_1, cout_29_2_1, cout_28_6_0, cout_28_7_0, cout_28_8_0);

wire sum_29_3_1, cout_29_3_1;

full_adder fa_29_3_1(sum_29_3_1, cout_29_3_1, cout_28_9_0, sum_29_0_0, sum_29_1_0);

wire sum_29_4_1, cout_29_4_1;

full_adder fa_29_4_1(sum_29_4_1, cout_29_4_1, sum_29_2_0, sum_29_3_0, sum_29_4_0);

wire sum_29_5_1, cout_29_5_1;

full_adder fa_29_5_1(sum_29_5_1, cout_29_5_1, sum_29_5_0, sum_29_6_0, sum_29_7_0);

wire sum_29_6_1, cout_29_6_1;

half_adder ha_29_6_1(sum_29_6_1, cout_29_6_1, sum_29_8_0, sum_29_9_0);

wire sum_30_0_1, cout_30_0_1;

full_adder fa_30_0_1(sum_30_0_1, cout_30_0_1, A0B30, cout_29_0_0, cout_29_1_0);

wire sum_30_1_1, cout_30_1_1;

full_adder fa_30_1_1(sum_30_1_1, cout_30_1_1, cout_29_2_0, cout_29_3_0, cout_29_4_0);

wire sum_30_2_1, cout_30_2_1;

full_adder fa_30_2_1(sum_30_2_1, cout_30_2_1, cout_29_5_0, cout_29_6_0, cout_29_7_0);

wire sum_30_3_1, cout_30_3_1;

full_adder fa_30_3_1(sum_30_3_1, cout_30_3_1, cout_29_8_0, cout_29_9_0, sum_30_0_0);

wire sum_30_4_1, cout_30_4_1;

full_adder fa_30_4_1(sum_30_4_1, cout_30_4_1, sum_30_1_0, sum_30_2_0, sum_30_3_0);

wire sum_30_5_1, cout_30_5_1;

full_adder fa_30_5_1(sum_30_5_1, cout_30_5_1, sum_30_4_0, sum_30_5_0, sum_30_6_0);

wire sum_30_6_1, cout_30_6_1;

full_adder fa_30_6_1(sum_30_6_1, cout_30_6_1, sum_30_7_0, sum_30_8_0, sum_30_9_0);

wire sum_31_0_1, cout_31_0_1;

full_adder fa_31_0_1(sum_31_0_1, cout_31_0_1, cout_30_0_0, cout_30_1_0, cout_30_2_0);

wire sum_31_1_1, cout_31_1_1;

full_adder fa_31_1_1(sum_31_1_1, cout_31_1_1, cout_30_3_0, cout_30_4_0, cout_30_5_0);

wire sum_31_2_1, cout_31_2_1;

full_adder fa_31_2_1(sum_31_2_1, cout_31_2_1, cout_30_6_0, cout_30_7_0, cout_30_8_0);

wire sum_31_3_1, cout_31_3_1;

full_adder fa_31_3_1(sum_31_3_1, cout_31_3_1, cout_30_9_0, sum_31_0_0, sum_31_1_0);

wire sum_31_4_1, cout_31_4_1;

full_adder fa_31_4_1(sum_31_4_1, cout_31_4_1, sum_31_2_0, sum_31_3_0, sum_31_4_0);

wire sum_31_5_1, cout_31_5_1;

full_adder fa_31_5_1(sum_31_5_1, cout_31_5_1, sum_31_5_0, sum_31_6_0, sum_31_7_0);

wire sum_31_6_1, cout_31_6_1;

full_adder fa_31_6_1(sum_31_6_1, cout_31_6_1, sum_31_8_0, sum_31_9_0, sum_31_10_0);

wire sum_32_0_1, cout_32_0_1;

full_adder fa_32_0_1(sum_32_0_1, cout_32_0_1, A1B31, cout_31_0_0, cout_31_1_0);

wire sum_32_1_1, cout_32_1_1;

full_adder fa_32_1_1(sum_32_1_1, cout_32_1_1, cout_31_2_0, cout_31_3_0, cout_31_4_0);

wire sum_32_2_1, cout_32_2_1;

full_adder fa_32_2_1(sum_32_2_1, cout_32_2_1, cout_31_5_0, cout_31_6_0, cout_31_7_0);

wire sum_32_3_1, cout_32_3_1;

full_adder fa_32_3_1(sum_32_3_1, cout_32_3_1, cout_31_8_0, cout_31_9_0, cout_31_10_0);

wire sum_32_4_1, cout_32_4_1;

full_adder fa_32_4_1(sum_32_4_1, cout_32_4_1, sum_32_0_0, sum_32_1_0, sum_32_2_0);

wire sum_32_5_1, cout_32_5_1;

full_adder fa_32_5_1(sum_32_5_1, cout_32_5_1, sum_32_3_0, sum_32_4_0, sum_32_5_0);

wire sum_32_6_1, cout_32_6_1;

full_adder fa_32_6_1(sum_32_6_1, cout_32_6_1, sum_32_6_0, sum_32_7_0, sum_32_8_0);

wire sum_33_0_1, cout_33_0_1;

full_adder fa_33_0_1(sum_33_0_1, cout_33_0_1, cout_32_0_0, cout_32_1_0, cout_32_2_0);

wire sum_33_1_1, cout_33_1_1;

full_adder fa_33_1_1(sum_33_1_1, cout_33_1_1, cout_32_3_0, cout_32_4_0, cout_32_5_0);

wire sum_33_2_1, cout_33_2_1;

full_adder fa_33_2_1(sum_33_2_1, cout_33_2_1, cout_32_6_0, cout_32_7_0, cout_32_8_0);

wire sum_33_3_1, cout_33_3_1;

full_adder fa_33_3_1(sum_33_3_1, cout_33_3_1, cout_32_9_0, sum_33_0_0, sum_33_1_0);

wire sum_33_4_1, cout_33_4_1;

full_adder fa_33_4_1(sum_33_4_1, cout_33_4_1, sum_33_2_0, sum_33_3_0, sum_33_4_0);

wire sum_33_5_1, cout_33_5_1;

full_adder fa_33_5_1(sum_33_5_1, cout_33_5_1, sum_33_5_0, sum_33_6_0, sum_33_7_0);

wire sum_33_6_1, cout_33_6_1;

half_adder ha_33_6_1(sum_33_6_1, cout_33_6_1, sum_33_8_0, sum_33_9_0);

wire sum_34_0_1, cout_34_0_1;

full_adder fa_34_0_1(sum_34_0_1, cout_34_0_1, cout_33_0_0, cout_33_1_0, cout_33_2_0);

wire sum_34_1_1, cout_34_1_1;

full_adder fa_34_1_1(sum_34_1_1, cout_34_1_1, cout_33_3_0, cout_33_4_0, cout_33_5_0);

wire sum_34_2_1, cout_34_2_1;

full_adder fa_34_2_1(sum_34_2_1, cout_34_2_1, cout_33_6_0, cout_33_7_0, cout_33_8_0);

wire sum_34_3_1, cout_34_3_1;

full_adder fa_34_3_1(sum_34_3_1, cout_34_3_1, cout_33_9_0, sum_34_0_0, sum_34_1_0);

wire sum_34_4_1, cout_34_4_1;

full_adder fa_34_4_1(sum_34_4_1, cout_34_4_1, sum_34_2_0, sum_34_3_0, sum_34_4_0);

wire sum_34_5_1, cout_34_5_1;

full_adder fa_34_5_1(sum_34_5_1, cout_34_5_1, sum_34_5_0, sum_34_6_0, sum_34_7_0);

wire sum_34_6_1, cout_34_6_1;

half_adder ha_34_6_1(sum_34_6_1, cout_34_6_1, sum_34_8_0, sum_34_9_0);

wire sum_35_0_1, cout_35_0_1;

full_adder fa_35_0_1(sum_35_0_1, cout_35_0_1, A4B31, cout_34_0_0, cout_34_1_0);

wire sum_35_1_1, cout_35_1_1;

full_adder fa_35_1_1(sum_35_1_1, cout_35_1_1, cout_34_2_0, cout_34_3_0, cout_34_4_0);

wire sum_35_2_1, cout_35_2_1;

full_adder fa_35_2_1(sum_35_2_1, cout_35_2_1, cout_34_5_0, cout_34_6_0, cout_34_7_0);

wire sum_35_3_1, cout_35_3_1;

full_adder fa_35_3_1(sum_35_3_1, cout_35_3_1, cout_34_8_0, cout_34_9_0, sum_35_0_0);

wire sum_35_4_1, cout_35_4_1;

full_adder fa_35_4_1(sum_35_4_1, cout_35_4_1, sum_35_1_0, sum_35_2_0, sum_35_3_0);

wire sum_35_5_1, cout_35_5_1;

full_adder fa_35_5_1(sum_35_5_1, cout_35_5_1, sum_35_4_0, sum_35_5_0, sum_35_6_0);

wire sum_35_6_1, cout_35_6_1;

half_adder ha_35_6_1(sum_35_6_1, cout_35_6_1, sum_35_7_0, sum_35_8_0);

wire sum_36_0_1, cout_36_0_1;

full_adder fa_36_0_1(sum_36_0_1, cout_36_0_1, cout_35_0_0, cout_35_1_0, cout_35_2_0);

wire sum_36_1_1, cout_36_1_1;

full_adder fa_36_1_1(sum_36_1_1, cout_36_1_1, cout_35_3_0, cout_35_4_0, cout_35_5_0);

wire sum_36_2_1, cout_36_2_1;

full_adder fa_36_2_1(sum_36_2_1, cout_36_2_1, cout_35_6_0, cout_35_7_0, cout_35_8_0);

wire sum_36_3_1, cout_36_3_1;

full_adder fa_36_3_1(sum_36_3_1, cout_36_3_1, sum_36_0_0, sum_36_1_0, sum_36_2_0);

wire sum_36_4_1, cout_36_4_1;

full_adder fa_36_4_1(sum_36_4_1, cout_36_4_1, sum_36_3_0, sum_36_4_0, sum_36_5_0);

wire sum_36_5_1, cout_36_5_1;

full_adder fa_36_5_1(sum_36_5_1, cout_36_5_1, sum_36_6_0, sum_36_7_0, sum_36_8_0);

wire sum_37_0_1, cout_37_0_1;

full_adder fa_37_0_1(sum_37_0_1, cout_37_0_1, cout_36_0_0, cout_36_1_0, cout_36_2_0);

wire sum_37_1_1, cout_37_1_1;

full_adder fa_37_1_1(sum_37_1_1, cout_37_1_1, cout_36_3_0, cout_36_4_0, cout_36_5_0);

wire sum_37_2_1, cout_37_2_1;

full_adder fa_37_2_1(sum_37_2_1, cout_37_2_1, cout_36_6_0, cout_36_7_0, cout_36_8_0);

wire sum_37_3_1, cout_37_3_1;

full_adder fa_37_3_1(sum_37_3_1, cout_37_3_1, sum_37_0_0, sum_37_1_0, sum_37_2_0);

wire sum_37_4_1, cout_37_4_1;

full_adder fa_37_4_1(sum_37_4_1, cout_37_4_1, sum_37_3_0, sum_37_4_0, sum_37_5_0);

wire sum_37_5_1, cout_37_5_1;

full_adder fa_37_5_1(sum_37_5_1, cout_37_5_1, sum_37_6_0, sum_37_7_0, sum_37_8_0);

wire sum_38_0_1, cout_38_0_1;

full_adder fa_38_0_1(sum_38_0_1, cout_38_0_1, A7B31, cout_37_0_0, cout_37_1_0);

wire sum_38_1_1, cout_38_1_1;

full_adder fa_38_1_1(sum_38_1_1, cout_38_1_1, cout_37_2_0, cout_37_3_0, cout_37_4_0);

wire sum_38_2_1, cout_38_2_1;

full_adder fa_38_2_1(sum_38_2_1, cout_38_2_1, cout_37_5_0, cout_37_6_0, cout_37_7_0);

wire sum_38_3_1, cout_38_3_1;

full_adder fa_38_3_1(sum_38_3_1, cout_38_3_1, cout_37_8_0, sum_38_0_0, sum_38_1_0);

wire sum_38_4_1, cout_38_4_1;

full_adder fa_38_4_1(sum_38_4_1, cout_38_4_1, sum_38_2_0, sum_38_3_0, sum_38_4_0);

wire sum_38_5_1, cout_38_5_1;

full_adder fa_38_5_1(sum_38_5_1, cout_38_5_1, sum_38_5_0, sum_38_6_0, sum_38_7_0);

wire sum_39_0_1, cout_39_0_1;

full_adder fa_39_0_1(sum_39_0_1, cout_39_0_1, cout_38_0_0, cout_38_1_0, cout_38_2_0);

wire sum_39_1_1, cout_39_1_1;

full_adder fa_39_1_1(sum_39_1_1, cout_39_1_1, cout_38_3_0, cout_38_4_0, cout_38_5_0);

wire sum_39_2_1, cout_39_2_1;

full_adder fa_39_2_1(sum_39_2_1, cout_39_2_1, cout_38_6_0, cout_38_7_0, sum_39_0_0);

wire sum_39_3_1, cout_39_3_1;

full_adder fa_39_3_1(sum_39_3_1, cout_39_3_1, sum_39_1_0, sum_39_2_0, sum_39_3_0);

wire sum_39_4_1, cout_39_4_1;

full_adder fa_39_4_1(sum_39_4_1, cout_39_4_1, sum_39_4_0, sum_39_5_0, sum_39_6_0);

wire sum_40_0_1, cout_40_0_1;

full_adder fa_40_0_1(sum_40_0_1, cout_40_0_1, cout_39_0_0, cout_39_1_0, cout_39_2_0);

wire sum_40_1_1, cout_40_1_1;

full_adder fa_40_1_1(sum_40_1_1, cout_40_1_1, cout_39_3_0, cout_39_4_0, cout_39_5_0);

wire sum_40_2_1, cout_40_2_1;

full_adder fa_40_2_1(sum_40_2_1, cout_40_2_1, cout_39_6_0, cout_39_7_0, sum_40_0_0);

wire sum_40_3_1, cout_40_3_1;

full_adder fa_40_3_1(sum_40_3_1, cout_40_3_1, sum_40_1_0, sum_40_2_0, sum_40_3_0);

wire sum_40_4_1, cout_40_4_1;

full_adder fa_40_4_1(sum_40_4_1, cout_40_4_1, sum_40_4_0, sum_40_5_0, sum_40_6_0);

wire sum_41_0_1, cout_41_0_1;

full_adder fa_41_0_1(sum_41_0_1, cout_41_0_1, A10B31, cout_40_0_0, cout_40_1_0);

wire sum_41_1_1, cout_41_1_1;

full_adder fa_41_1_1(sum_41_1_1, cout_41_1_1, cout_40_2_0, cout_40_3_0, cout_40_4_0);

wire sum_41_2_1, cout_41_2_1;

full_adder fa_41_2_1(sum_41_2_1, cout_41_2_1, cout_40_5_0, cout_40_6_0, cout_40_7_0);

wire sum_41_3_1, cout_41_3_1;

full_adder fa_41_3_1(sum_41_3_1, cout_41_3_1, sum_41_0_0, sum_41_1_0, sum_41_2_0);

wire sum_41_4_1, cout_41_4_1;

full_adder fa_41_4_1(sum_41_4_1, cout_41_4_1, sum_41_3_0, sum_41_4_0, sum_41_5_0);

wire sum_42_0_1, cout_42_0_1;

full_adder fa_42_0_1(sum_42_0_1, cout_42_0_1, cout_41_0_0, cout_41_1_0, cout_41_2_0);

wire sum_42_1_1, cout_42_1_1;

full_adder fa_42_1_1(sum_42_1_1, cout_42_1_1, cout_41_3_0, cout_41_4_0, cout_41_5_0);

wire sum_42_2_1, cout_42_2_1;

full_adder fa_42_2_1(sum_42_2_1, cout_42_2_1, cout_41_6_0, sum_42_0_0, sum_42_1_0);

wire sum_42_3_1, cout_42_3_1;

full_adder fa_42_3_1(sum_42_3_1, cout_42_3_1, sum_42_2_0, sum_42_3_0, sum_42_4_0);

wire sum_42_4_1, cout_42_4_1;

half_adder ha_42_4_1(sum_42_4_1, cout_42_4_1, sum_42_5_0, sum_42_6_0);

wire sum_43_0_1, cout_43_0_1;

full_adder fa_43_0_1(sum_43_0_1, cout_43_0_1, cout_42_0_0, cout_42_1_0, cout_42_2_0);

wire sum_43_1_1, cout_43_1_1;

full_adder fa_43_1_1(sum_43_1_1, cout_43_1_1, cout_42_3_0, cout_42_4_0, cout_42_5_0);

wire sum_43_2_1, cout_43_2_1;

full_adder fa_43_2_1(sum_43_2_1, cout_43_2_1, cout_42_6_0, sum_43_0_0, sum_43_1_0);

wire sum_43_3_1, cout_43_3_1;

full_adder fa_43_3_1(sum_43_3_1, cout_43_3_1, sum_43_2_0, sum_43_3_0, sum_43_4_0);

wire sum_43_4_1, cout_43_4_1;

half_adder ha_43_4_1(sum_43_4_1, cout_43_4_1, sum_43_5_0, sum_43_6_0);

wire sum_44_0_1, cout_44_0_1;

full_adder fa_44_0_1(sum_44_0_1, cout_44_0_1, A13B31, cout_43_0_0, cout_43_1_0);

wire sum_44_1_1, cout_44_1_1;

full_adder fa_44_1_1(sum_44_1_1, cout_44_1_1, cout_43_2_0, cout_43_3_0, cout_43_4_0);

wire sum_44_2_1, cout_44_2_1;

full_adder fa_44_2_1(sum_44_2_1, cout_44_2_1, cout_43_5_0, cout_43_6_0, sum_44_0_0);

wire sum_44_3_1, cout_44_3_1;

full_adder fa_44_3_1(sum_44_3_1, cout_44_3_1, sum_44_1_0, sum_44_2_0, sum_44_3_0);

wire sum_44_4_1, cout_44_4_1;

half_adder ha_44_4_1(sum_44_4_1, cout_44_4_1, sum_44_4_0, sum_44_5_0);

wire sum_45_0_1, cout_45_0_1;

full_adder fa_45_0_1(sum_45_0_1, cout_45_0_1, cout_44_0_0, cout_44_1_0, cout_44_2_0);

wire sum_45_1_1, cout_45_1_1;

full_adder fa_45_1_1(sum_45_1_1, cout_45_1_1, cout_44_3_0, cout_44_4_0, cout_44_5_0);

wire sum_45_2_1, cout_45_2_1;

full_adder fa_45_2_1(sum_45_2_1, cout_45_2_1, sum_45_0_0, sum_45_1_0, sum_45_2_0);

wire sum_45_3_1, cout_45_3_1;

full_adder fa_45_3_1(sum_45_3_1, cout_45_3_1, sum_45_3_0, sum_45_4_0, sum_45_5_0);

wire sum_46_0_1, cout_46_0_1;

full_adder fa_46_0_1(sum_46_0_1, cout_46_0_1, cout_45_0_0, cout_45_1_0, cout_45_2_0);

wire sum_46_1_1, cout_46_1_1;

full_adder fa_46_1_1(sum_46_1_1, cout_46_1_1, cout_45_3_0, cout_45_4_0, cout_45_5_0);

wire sum_46_2_1, cout_46_2_1;

full_adder fa_46_2_1(sum_46_2_1, cout_46_2_1, sum_46_0_0, sum_46_1_0, sum_46_2_0);

wire sum_46_3_1, cout_46_3_1;

full_adder fa_46_3_1(sum_46_3_1, cout_46_3_1, sum_46_3_0, sum_46_4_0, sum_46_5_0);

wire sum_47_0_1, cout_47_0_1;

full_adder fa_47_0_1(sum_47_0_1, cout_47_0_1, A16B31, cout_46_0_0, cout_46_1_0);

wire sum_47_1_1, cout_47_1_1;

full_adder fa_47_1_1(sum_47_1_1, cout_47_1_1, cout_46_2_0, cout_46_3_0, cout_46_4_0);

wire sum_47_2_1, cout_47_2_1;

full_adder fa_47_2_1(sum_47_2_1, cout_47_2_1, cout_46_5_0, sum_47_0_0, sum_47_1_0);

wire sum_47_3_1, cout_47_3_1;

full_adder fa_47_3_1(sum_47_3_1, cout_47_3_1, sum_47_2_0, sum_47_3_0, sum_47_4_0);

wire sum_48_0_1, cout_48_0_1;

full_adder fa_48_0_1(sum_48_0_1, cout_48_0_1, cout_47_0_0, cout_47_1_0, cout_47_2_0);

wire sum_48_1_1, cout_48_1_1;

full_adder fa_48_1_1(sum_48_1_1, cout_48_1_1, cout_47_3_0, cout_47_4_0, sum_48_0_0);

wire sum_48_2_1, cout_48_2_1;

full_adder fa_48_2_1(sum_48_2_1, cout_48_2_1, sum_48_1_0, sum_48_2_0, sum_48_3_0);

wire sum_49_0_1, cout_49_0_1;

full_adder fa_49_0_1(sum_49_0_1, cout_49_0_1, cout_48_0_0, cout_48_1_0, cout_48_2_0);

wire sum_49_1_1, cout_49_1_1;

full_adder fa_49_1_1(sum_49_1_1, cout_49_1_1, cout_48_3_0, cout_48_4_0, sum_49_0_0);

wire sum_49_2_1, cout_49_2_1;

full_adder fa_49_2_1(sum_49_2_1, cout_49_2_1, sum_49_1_0, sum_49_2_0, sum_49_3_0);

wire sum_50_0_1, cout_50_0_1;

full_adder fa_50_0_1(sum_50_0_1, cout_50_0_1, A19B31, cout_49_0_0, cout_49_1_0);

wire sum_50_1_1, cout_50_1_1;

full_adder fa_50_1_1(sum_50_1_1, cout_50_1_1, cout_49_2_0, cout_49_3_0, cout_49_4_0);

wire sum_50_2_1, cout_50_2_1;

full_adder fa_50_2_1(sum_50_2_1, cout_50_2_1, sum_50_0_0, sum_50_1_0, sum_50_2_0);

wire sum_51_0_1, cout_51_0_1;

full_adder fa_51_0_1(sum_51_0_1, cout_51_0_1, cout_50_0_0, cout_50_1_0, cout_50_2_0);

wire sum_51_1_1, cout_51_1_1;

full_adder fa_51_1_1(sum_51_1_1, cout_51_1_1, cout_50_3_0, sum_51_0_0, sum_51_1_0);

wire sum_51_2_1, cout_51_2_1;

half_adder ha_51_2_1(sum_51_2_1, cout_51_2_1, sum_51_2_0, sum_51_3_0);

wire sum_52_0_1, cout_52_0_1;

full_adder fa_52_0_1(sum_52_0_1, cout_52_0_1, cout_51_0_0, cout_51_1_0, cout_51_2_0);

wire sum_52_1_1, cout_52_1_1;

full_adder fa_52_1_1(sum_52_1_1, cout_52_1_1, cout_51_3_0, sum_52_0_0, sum_52_1_0);

wire sum_52_2_1, cout_52_2_1;

half_adder ha_52_2_1(sum_52_2_1, cout_52_2_1, sum_52_2_0, sum_52_3_0);

wire sum_53_0_1, cout_53_0_1;

full_adder fa_53_0_1(sum_53_0_1, cout_53_0_1, A22B31, cout_52_0_0, cout_52_1_0);

wire sum_53_1_1, cout_53_1_1;

full_adder fa_53_1_1(sum_53_1_1, cout_53_1_1, cout_52_2_0, cout_52_3_0, sum_53_0_0);

wire sum_53_2_1, cout_53_2_1;

half_adder ha_53_2_1(sum_53_2_1, cout_53_2_1, sum_53_1_0, sum_53_2_0);

wire sum_54_0_1, cout_54_0_1;

full_adder fa_54_0_1(sum_54_0_1, cout_54_0_1, cout_53_0_0, cout_53_1_0, cout_53_2_0);

wire sum_54_1_1, cout_54_1_1;

full_adder fa_54_1_1(sum_54_1_1, cout_54_1_1, sum_54_0_0, sum_54_1_0, sum_54_2_0);

wire sum_55_0_1, cout_55_0_1;

full_adder fa_55_0_1(sum_55_0_1, cout_55_0_1, cout_54_0_0, cout_54_1_0, cout_54_2_0);

wire sum_55_1_1, cout_55_1_1;

full_adder fa_55_1_1(sum_55_1_1, cout_55_1_1, sum_55_0_0, sum_55_1_0, sum_55_2_0);

wire sum_56_0_1, cout_56_0_1;

full_adder fa_56_0_1(sum_56_0_1, cout_56_0_1, A25B31, cout_55_0_0, cout_55_1_0);

wire sum_56_1_1, cout_56_1_1;

full_adder fa_56_1_1(sum_56_1_1, cout_56_1_1, cout_55_2_0, sum_56_0_0, sum_56_1_0);

wire sum_57_0_1, cout_57_0_1;

full_adder fa_57_0_1(sum_57_0_1, cout_57_0_1, cout_56_0_0, cout_56_1_0, sum_57_0_0);

wire sum_58_0_1, cout_58_0_1;

full_adder fa_58_0_1(sum_58_0_1, cout_58_0_1, cout_57_0_0, cout_57_1_0, sum_58_0_0);

wire sum_59_0_1, cout_59_0_1;

full_adder fa_59_0_1(sum_59_0_1, cout_59_0_1, A28B31, cout_58_0_0, cout_58_1_0);

wire sum_5_0_2, cout_5_0_2;

half_adder ha_5_0_2(sum_5_0_2, cout_5_0_2, sum_5_1_0, cout_4_0_1);

wire sum_6_0_2, cout_6_0_2;

full_adder fa_6_0_2(sum_6_0_2, cout_6_0_2, cout_5_0_1, sum_6_0_1, sum_6_1_1);

wire sum_7_0_2, cout_7_0_2;

full_adder fa_7_0_2(sum_7_0_2, cout_7_0_2, cout_6_0_1, cout_6_1_1, sum_7_0_1);

wire sum_8_0_2, cout_8_0_2;

full_adder fa_8_0_2(sum_8_0_2, cout_8_0_2, cout_7_0_1, cout_7_1_1, sum_8_0_1);

wire sum_9_0_2, cout_9_0_2;

full_adder fa_9_0_2(sum_9_0_2, cout_9_0_2, sum_9_2_0, cout_8_0_1, cout_8_1_1);

wire sum_9_1_2, cout_9_1_2;

half_adder ha_9_1_2(sum_9_1_2, cout_9_1_2, sum_9_0_1, sum_9_1_1);

wire sum_10_0_2, cout_10_0_2;

full_adder fa_10_0_2(sum_10_0_2, cout_10_0_2, sum_10_3_0, cout_9_0_1, cout_9_1_1);

wire sum_10_1_2, cout_10_1_2;

half_adder ha_10_1_2(sum_10_1_2, cout_10_1_2, sum_10_0_1, sum_10_1_1);

wire sum_11_0_2, cout_11_0_2;

full_adder fa_11_0_2(sum_11_0_2, cout_11_0_2, cout_10_0_1, cout_10_1_1, sum_11_0_1);

wire sum_11_1_2, cout_11_1_2;

half_adder ha_11_1_2(sum_11_1_2, cout_11_1_2, sum_11_1_1, sum_11_2_1);

wire sum_12_0_2, cout_12_0_2;

full_adder fa_12_0_2(sum_12_0_2, cout_12_0_2, cout_11_0_1, cout_11_1_1, cout_11_2_1);

wire sum_12_1_2, cout_12_1_2;

full_adder fa_12_1_2(sum_12_1_2, cout_12_1_2, sum_12_0_1, sum_12_1_1, sum_12_2_1);

wire sum_13_0_2, cout_13_0_2;

full_adder fa_13_0_2(sum_13_0_2, cout_13_0_2, cout_12_0_1, cout_12_1_1, cout_12_2_1);

wire sum_13_1_2, cout_13_1_2;

full_adder fa_13_1_2(sum_13_1_2, cout_13_1_2, sum_13_0_1, sum_13_1_1, sum_13_2_1);

wire sum_14_0_2, cout_14_0_2;

full_adder fa_14_0_2(sum_14_0_2, cout_14_0_2, sum_14_4_0, cout_13_0_1, cout_13_1_1);

wire sum_14_1_2, cout_14_1_2;

full_adder fa_14_1_2(sum_14_1_2, cout_14_1_2, cout_13_2_1, sum_14_0_1, sum_14_1_1);

wire sum_15_0_2, cout_15_0_2;

full_adder fa_15_0_2(sum_15_0_2, cout_15_0_2, cout_14_0_1, cout_14_1_1, cout_14_2_1);

wire sum_15_1_2, cout_15_1_2;

full_adder fa_15_1_2(sum_15_1_2, cout_15_1_2, sum_15_0_1, sum_15_1_1, sum_15_2_1);

wire sum_16_0_2, cout_16_0_2;

full_adder fa_16_0_2(sum_16_0_2, cout_16_0_2, cout_15_0_1, cout_15_1_1, cout_15_2_1);

wire sum_16_1_2, cout_16_1_2;

full_adder fa_16_1_2(sum_16_1_2, cout_16_1_2, cout_15_3_1, sum_16_0_1, sum_16_1_1);

wire sum_16_2_2, cout_16_2_2;

half_adder ha_16_2_2(sum_16_2_2, cout_16_2_2, sum_16_2_1, sum_16_3_1);

wire sum_17_0_2, cout_17_0_2;

full_adder fa_17_0_2(sum_17_0_2, cout_17_0_2, cout_16_0_1, cout_16_1_1, cout_16_2_1);

wire sum_17_1_2, cout_17_1_2;

full_adder fa_17_1_2(sum_17_1_2, cout_17_1_2, cout_16_3_1, sum_17_0_1, sum_17_1_1);

wire sum_17_2_2, cout_17_2_2;

half_adder ha_17_2_2(sum_17_2_2, cout_17_2_2, sum_17_2_1, sum_17_3_1);

wire sum_18_0_2, cout_18_0_2;

full_adder fa_18_0_2(sum_18_0_2, cout_18_0_2, sum_18_5_0, cout_17_0_1, cout_17_1_1);

wire sum_18_1_2, cout_18_1_2;

full_adder fa_18_1_2(sum_18_1_2, cout_18_1_2, cout_17_2_1, cout_17_3_1, sum_18_0_1);

wire sum_18_2_2, cout_18_2_2;

full_adder fa_18_2_2(sum_18_2_2, cout_18_2_2, sum_18_1_1, sum_18_2_1, sum_18_3_1);

wire sum_19_0_2, cout_19_0_2;

full_adder fa_19_0_2(sum_19_0_2, cout_19_0_2, sum_19_6_0, cout_18_0_1, cout_18_1_1);

wire sum_19_1_2, cout_19_1_2;

full_adder fa_19_1_2(sum_19_1_2, cout_19_1_2, cout_18_2_1, cout_18_3_1, sum_19_0_1);

wire sum_19_2_2, cout_19_2_2;

full_adder fa_19_2_2(sum_19_2_2, cout_19_2_2, sum_19_1_1, sum_19_2_1, sum_19_3_1);

wire sum_20_0_2, cout_20_0_2;

full_adder fa_20_0_2(sum_20_0_2, cout_20_0_2, cout_19_0_1, cout_19_1_1, cout_19_2_1);

wire sum_20_1_2, cout_20_1_2;

full_adder fa_20_1_2(sum_20_1_2, cout_20_1_2, cout_19_3_1, sum_20_0_1, sum_20_1_1);

wire sum_20_2_2, cout_20_2_2;

full_adder fa_20_2_2(sum_20_2_2, cout_20_2_2, sum_20_2_1, sum_20_3_1, sum_20_4_1);

wire sum_21_0_2, cout_21_0_2;

full_adder fa_21_0_2(sum_21_0_2, cout_21_0_2, cout_20_0_1, cout_20_1_1, cout_20_2_1);

wire sum_21_1_2, cout_21_1_2;

full_adder fa_21_1_2(sum_21_1_2, cout_21_1_2, cout_20_3_1, cout_20_4_1, sum_21_0_1);

wire sum_21_2_2, cout_21_2_2;

full_adder fa_21_2_2(sum_21_2_2, cout_21_2_2, sum_21_1_1, sum_21_2_1, sum_21_3_1);

wire sum_22_0_2, cout_22_0_2;

full_adder fa_22_0_2(sum_22_0_2, cout_22_0_2, cout_21_0_1, cout_21_1_1, cout_21_2_1);

wire sum_22_1_2, cout_22_1_2;

full_adder fa_22_1_2(sum_22_1_2, cout_22_1_2, cout_21_3_1, cout_21_4_1, sum_22_0_1);

wire sum_22_2_2, cout_22_2_2;

full_adder fa_22_2_2(sum_22_2_2, cout_22_2_2, sum_22_1_1, sum_22_2_1, sum_22_3_1);

wire sum_23_0_2, cout_23_0_2;

full_adder fa_23_0_2(sum_23_0_2, cout_23_0_2, sum_23_7_0, cout_22_0_1, cout_22_1_1);

wire sum_23_1_2, cout_23_1_2;

full_adder fa_23_1_2(sum_23_1_2, cout_23_1_2, cout_22_2_1, cout_22_3_1, cout_22_4_1);

wire sum_23_2_2, cout_23_2_2;

full_adder fa_23_2_2(sum_23_2_2, cout_23_2_2, sum_23_0_1, sum_23_1_1, sum_23_2_1);

wire sum_23_3_2, cout_23_3_2;

half_adder ha_23_3_2(sum_23_3_2, cout_23_3_2, sum_23_3_1, sum_23_4_1);

wire sum_24_0_2, cout_24_0_2;

full_adder fa_24_0_2(sum_24_0_2, cout_24_0_2, cout_23_0_1, cout_23_1_1, cout_23_2_1);

wire sum_24_1_2, cout_24_1_2;

full_adder fa_24_1_2(sum_24_1_2, cout_24_1_2, cout_23_3_1, cout_23_4_1, sum_24_0_1);

wire sum_24_2_2, cout_24_2_2;

full_adder fa_24_2_2(sum_24_2_2, cout_24_2_2, sum_24_1_1, sum_24_2_1, sum_24_3_1);

wire sum_24_3_2, cout_24_3_2;

half_adder ha_24_3_2(sum_24_3_2, cout_24_3_2, sum_24_4_1, sum_24_5_1);

wire sum_25_0_2, cout_25_0_2;

full_adder fa_25_0_2(sum_25_0_2, cout_25_0_2, cout_24_0_1, cout_24_1_1, cout_24_2_1);

wire sum_25_1_2, cout_25_1_2;

full_adder fa_25_1_2(sum_25_1_2, cout_25_1_2, cout_24_3_1, cout_24_4_1, cout_24_5_1);

wire sum_25_2_2, cout_25_2_2;

full_adder fa_25_2_2(sum_25_2_2, cout_25_2_2, sum_25_0_1, sum_25_1_1, sum_25_2_1);

wire sum_25_3_2, cout_25_3_2;

full_adder fa_25_3_2(sum_25_3_2, cout_25_3_2, sum_25_3_1, sum_25_4_1, sum_25_5_1);

wire sum_26_0_2, cout_26_0_2;

full_adder fa_26_0_2(sum_26_0_2, cout_26_0_2, cout_25_0_1, cout_25_1_1, cout_25_2_1);

wire sum_26_1_2, cout_26_1_2;

full_adder fa_26_1_2(sum_26_1_2, cout_26_1_2, cout_25_3_1, cout_25_4_1, cout_25_5_1);

wire sum_26_2_2, cout_26_2_2;

full_adder fa_26_2_2(sum_26_2_2, cout_26_2_2, sum_26_0_1, sum_26_1_1, sum_26_2_1);

wire sum_26_3_2, cout_26_3_2;

full_adder fa_26_3_2(sum_26_3_2, cout_26_3_2, sum_26_3_1, sum_26_4_1, sum_26_5_1);

wire sum_27_0_2, cout_27_0_2;

full_adder fa_27_0_2(sum_27_0_2, cout_27_0_2, sum_27_8_0, cout_26_0_1, cout_26_1_1);

wire sum_27_1_2, cout_27_1_2;

full_adder fa_27_1_2(sum_27_1_2, cout_27_1_2, cout_26_2_1, cout_26_3_1, cout_26_4_1);

wire sum_27_2_2, cout_27_2_2;

full_adder fa_27_2_2(sum_27_2_2, cout_27_2_2, cout_26_5_1, sum_27_0_1, sum_27_1_1);

wire sum_27_3_2, cout_27_3_2;

full_adder fa_27_3_2(sum_27_3_2, cout_27_3_2, sum_27_2_1, sum_27_3_1, sum_27_4_1);

wire sum_28_0_2, cout_28_0_2;

full_adder fa_28_0_2(sum_28_0_2, cout_28_0_2, sum_28_9_0, cout_27_0_1, cout_27_1_1);

wire sum_28_1_2, cout_28_1_2;

full_adder fa_28_1_2(sum_28_1_2, cout_28_1_2, cout_27_2_1, cout_27_3_1, cout_27_4_1);

wire sum_28_2_2, cout_28_2_2;

full_adder fa_28_2_2(sum_28_2_2, cout_28_2_2, cout_27_5_1, sum_28_0_1, sum_28_1_1);

wire sum_28_3_2, cout_28_3_2;

full_adder fa_28_3_2(sum_28_3_2, cout_28_3_2, sum_28_2_1, sum_28_3_1, sum_28_4_1);

wire sum_29_0_2, cout_29_0_2;

full_adder fa_29_0_2(sum_29_0_2, cout_29_0_2, cout_28_0_1, cout_28_1_1, cout_28_2_1);

wire sum_29_1_2, cout_29_1_2;

full_adder fa_29_1_2(sum_29_1_2, cout_29_1_2, cout_28_3_1, cout_28_4_1, cout_28_5_1);

wire sum_29_2_2, cout_29_2_2;

full_adder fa_29_2_2(sum_29_2_2, cout_29_2_2, sum_29_0_1, sum_29_1_1, sum_29_2_1);

wire sum_29_3_2, cout_29_3_2;

full_adder fa_29_3_2(sum_29_3_2, cout_29_3_2, sum_29_3_1, sum_29_4_1, sum_29_5_1);

wire sum_30_0_2, cout_30_0_2;

full_adder fa_30_0_2(sum_30_0_2, cout_30_0_2, cout_29_0_1, cout_29_1_1, cout_29_2_1);

wire sum_30_1_2, cout_30_1_2;

full_adder fa_30_1_2(sum_30_1_2, cout_30_1_2, cout_29_3_1, cout_29_4_1, cout_29_5_1);

wire sum_30_2_2, cout_30_2_2;

full_adder fa_30_2_2(sum_30_2_2, cout_30_2_2, cout_29_6_1, sum_30_0_1, sum_30_1_1);

wire sum_30_3_2, cout_30_3_2;

full_adder fa_30_3_2(sum_30_3_2, cout_30_3_2, sum_30_2_1, sum_30_3_1, sum_30_4_1);

wire sum_30_4_2, cout_30_4_2;

half_adder ha_30_4_2(sum_30_4_2, cout_30_4_2, sum_30_5_1, sum_30_6_1);

wire sum_31_0_2, cout_31_0_2;

full_adder fa_31_0_2(sum_31_0_2, cout_31_0_2, cout_30_0_1, cout_30_1_1, cout_30_2_1);

wire sum_31_1_2, cout_31_1_2;

full_adder fa_31_1_2(sum_31_1_2, cout_31_1_2, cout_30_3_1, cout_30_4_1, cout_30_5_1);

wire sum_31_2_2, cout_31_2_2;

full_adder fa_31_2_2(sum_31_2_2, cout_31_2_2, cout_30_6_1, sum_31_0_1, sum_31_1_1);

wire sum_31_3_2, cout_31_3_2;

full_adder fa_31_3_2(sum_31_3_2, cout_31_3_2, sum_31_2_1, sum_31_3_1, sum_31_4_1);

wire sum_31_4_2, cout_31_4_2;

half_adder ha_31_4_2(sum_31_4_2, cout_31_4_2, sum_31_5_1, sum_31_6_1);

wire sum_32_0_2, cout_32_0_2;

full_adder fa_32_0_2(sum_32_0_2, cout_32_0_2, sum_32_9_0, cout_31_0_1, cout_31_1_1);

wire sum_32_1_2, cout_32_1_2;

full_adder fa_32_1_2(sum_32_1_2, cout_32_1_2, cout_31_2_1, cout_31_3_1, cout_31_4_1);

wire sum_32_2_2, cout_32_2_2;

full_adder fa_32_2_2(sum_32_2_2, cout_32_2_2, cout_31_5_1, cout_31_6_1, sum_32_0_1);

wire sum_32_3_2, cout_32_3_2;

full_adder fa_32_3_2(sum_32_3_2, cout_32_3_2, sum_32_1_1, sum_32_2_1, sum_32_3_1);

wire sum_32_4_2, cout_32_4_2;

full_adder fa_32_4_2(sum_32_4_2, cout_32_4_2, sum_32_4_1, sum_32_5_1, sum_32_6_1);

wire sum_33_0_2, cout_33_0_2;

full_adder fa_33_0_2(sum_33_0_2, cout_33_0_2, cout_32_0_1, cout_32_1_1, cout_32_2_1);

wire sum_33_1_2, cout_33_1_2;

full_adder fa_33_1_2(sum_33_1_2, cout_33_1_2, cout_32_3_1, cout_32_4_1, cout_32_5_1);

wire sum_33_2_2, cout_33_2_2;

full_adder fa_33_2_2(sum_33_2_2, cout_33_2_2, cout_32_6_1, sum_33_0_1, sum_33_1_1);

wire sum_33_3_2, cout_33_3_2;

full_adder fa_33_3_2(sum_33_3_2, cout_33_3_2, sum_33_2_1, sum_33_3_1, sum_33_4_1);

wire sum_33_4_2, cout_33_4_2;

half_adder ha_33_4_2(sum_33_4_2, cout_33_4_2, sum_33_5_1, sum_33_6_1);

wire sum_34_0_2, cout_34_0_2;

full_adder fa_34_0_2(sum_34_0_2, cout_34_0_2, cout_33_0_1, cout_33_1_1, cout_33_2_1);

wire sum_34_1_2, cout_34_1_2;

full_adder fa_34_1_2(sum_34_1_2, cout_34_1_2, cout_33_3_1, cout_33_4_1, cout_33_5_1);

wire sum_34_2_2, cout_34_2_2;

full_adder fa_34_2_2(sum_34_2_2, cout_34_2_2, cout_33_6_1, sum_34_0_1, sum_34_1_1);

wire sum_34_3_2, cout_34_3_2;

full_adder fa_34_3_2(sum_34_3_2, cout_34_3_2, sum_34_2_1, sum_34_3_1, sum_34_4_1);

wire sum_34_4_2, cout_34_4_2;

half_adder ha_34_4_2(sum_34_4_2, cout_34_4_2, sum_34_5_1, sum_34_6_1);

wire sum_35_0_2, cout_35_0_2;

full_adder fa_35_0_2(sum_35_0_2, cout_35_0_2, cout_34_0_1, cout_34_1_1, cout_34_2_1);

wire sum_35_1_2, cout_35_1_2;

full_adder fa_35_1_2(sum_35_1_2, cout_35_1_2, cout_34_3_1, cout_34_4_1, cout_34_5_1);

wire sum_35_2_2, cout_35_2_2;

full_adder fa_35_2_2(sum_35_2_2, cout_35_2_2, cout_34_6_1, sum_35_0_1, sum_35_1_1);

wire sum_35_3_2, cout_35_3_2;

full_adder fa_35_3_2(sum_35_3_2, cout_35_3_2, sum_35_2_1, sum_35_3_1, sum_35_4_1);

wire sum_35_4_2, cout_35_4_2;

half_adder ha_35_4_2(sum_35_4_2, cout_35_4_2, sum_35_5_1, sum_35_6_1);

wire sum_36_0_2, cout_36_0_2;

full_adder fa_36_0_2(sum_36_0_2, cout_36_0_2, cout_35_0_1, cout_35_1_1, cout_35_2_1);

wire sum_36_1_2, cout_36_1_2;

full_adder fa_36_1_2(sum_36_1_2, cout_36_1_2, cout_35_3_1, cout_35_4_1, cout_35_5_1);

wire sum_36_2_2, cout_36_2_2;

full_adder fa_36_2_2(sum_36_2_2, cout_36_2_2, cout_35_6_1, sum_36_0_1, sum_36_1_1);

wire sum_36_3_2, cout_36_3_2;

full_adder fa_36_3_2(sum_36_3_2, cout_36_3_2, sum_36_2_1, sum_36_3_1, sum_36_4_1);

wire sum_37_0_2, cout_37_0_2;

full_adder fa_37_0_2(sum_37_0_2, cout_37_0_2, cout_36_0_1, cout_36_1_1, cout_36_2_1);

wire sum_37_1_2, cout_37_1_2;

full_adder fa_37_1_2(sum_37_1_2, cout_37_1_2, cout_36_3_1, cout_36_4_1, cout_36_5_1);

wire sum_37_2_2, cout_37_2_2;

full_adder fa_37_2_2(sum_37_2_2, cout_37_2_2, sum_37_0_1, sum_37_1_1, sum_37_2_1);

wire sum_37_3_2, cout_37_3_2;

full_adder fa_37_3_2(sum_37_3_2, cout_37_3_2, sum_37_3_1, sum_37_4_1, sum_37_5_1);

wire sum_38_0_2, cout_38_0_2;

full_adder fa_38_0_2(sum_38_0_2, cout_38_0_2, cout_37_0_1, cout_37_1_1, cout_37_2_1);

wire sum_38_1_2, cout_38_1_2;

full_adder fa_38_1_2(sum_38_1_2, cout_38_1_2, cout_37_3_1, cout_37_4_1, cout_37_5_1);

wire sum_38_2_2, cout_38_2_2;

full_adder fa_38_2_2(sum_38_2_2, cout_38_2_2, sum_38_0_1, sum_38_1_1, sum_38_2_1);

wire sum_38_3_2, cout_38_3_2;

full_adder fa_38_3_2(sum_38_3_2, cout_38_3_2, sum_38_3_1, sum_38_4_1, sum_38_5_1);

wire sum_39_0_2, cout_39_0_2;

full_adder fa_39_0_2(sum_39_0_2, cout_39_0_2, sum_39_7_0, cout_38_0_1, cout_38_1_1);

wire sum_39_1_2, cout_39_1_2;

full_adder fa_39_1_2(sum_39_1_2, cout_39_1_2, cout_38_2_1, cout_38_3_1, cout_38_4_1);

wire sum_39_2_2, cout_39_2_2;

full_adder fa_39_2_2(sum_39_2_2, cout_39_2_2, cout_38_5_1, sum_39_0_1, sum_39_1_1);

wire sum_39_3_2, cout_39_3_2;

full_adder fa_39_3_2(sum_39_3_2, cout_39_3_2, sum_39_2_1, sum_39_3_1, sum_39_4_1);

wire sum_40_0_2, cout_40_0_2;

full_adder fa_40_0_2(sum_40_0_2, cout_40_0_2, sum_40_7_0, cout_39_0_1, cout_39_1_1);

wire sum_40_1_2, cout_40_1_2;

full_adder fa_40_1_2(sum_40_1_2, cout_40_1_2, cout_39_2_1, cout_39_3_1, cout_39_4_1);

wire sum_40_2_2, cout_40_2_2;

full_adder fa_40_2_2(sum_40_2_2, cout_40_2_2, sum_40_0_1, sum_40_1_1, sum_40_2_1);

wire sum_40_3_2, cout_40_3_2;

half_adder ha_40_3_2(sum_40_3_2, cout_40_3_2, sum_40_3_1, sum_40_4_1);

wire sum_41_0_2, cout_41_0_2;

full_adder fa_41_0_2(sum_41_0_2, cout_41_0_2, sum_41_6_0, cout_40_0_1, cout_40_1_1);

wire sum_41_1_2, cout_41_1_2;

full_adder fa_41_1_2(sum_41_1_2, cout_41_1_2, cout_40_2_1, cout_40_3_1, cout_40_4_1);

wire sum_41_2_2, cout_41_2_2;

full_adder fa_41_2_2(sum_41_2_2, cout_41_2_2, sum_41_0_1, sum_41_1_1, sum_41_2_1);

wire sum_41_3_2, cout_41_3_2;

half_adder ha_41_3_2(sum_41_3_2, cout_41_3_2, sum_41_3_1, sum_41_4_1);

wire sum_42_0_2, cout_42_0_2;

full_adder fa_42_0_2(sum_42_0_2, cout_42_0_2, cout_41_0_1, cout_41_1_1, cout_41_2_1);

wire sum_42_1_2, cout_42_1_2;

full_adder fa_42_1_2(sum_42_1_2, cout_42_1_2, cout_41_3_1, cout_41_4_1, sum_42_0_1);

wire sum_42_2_2, cout_42_2_2;

full_adder fa_42_2_2(sum_42_2_2, cout_42_2_2, sum_42_1_1, sum_42_2_1, sum_42_3_1);

wire sum_43_0_2, cout_43_0_2;

full_adder fa_43_0_2(sum_43_0_2, cout_43_0_2, cout_42_0_1, cout_42_1_1, cout_42_2_1);

wire sum_43_1_2, cout_43_1_2;

full_adder fa_43_1_2(sum_43_1_2, cout_43_1_2, cout_42_3_1, cout_42_4_1, sum_43_0_1);

wire sum_43_2_2, cout_43_2_2;

full_adder fa_43_2_2(sum_43_2_2, cout_43_2_2, sum_43_1_1, sum_43_2_1, sum_43_3_1);

wire sum_44_0_2, cout_44_0_2;

full_adder fa_44_0_2(sum_44_0_2, cout_44_0_2, cout_43_0_1, cout_43_1_1, cout_43_2_1);

wire sum_44_1_2, cout_44_1_2;

full_adder fa_44_1_2(sum_44_1_2, cout_44_1_2, cout_43_3_1, cout_43_4_1, sum_44_0_1);

wire sum_44_2_2, cout_44_2_2;

full_adder fa_44_2_2(sum_44_2_2, cout_44_2_2, sum_44_1_1, sum_44_2_1, sum_44_3_1);

wire sum_45_0_2, cout_45_0_2;

full_adder fa_45_0_2(sum_45_0_2, cout_45_0_2, cout_44_0_1, cout_44_1_1, cout_44_2_1);

wire sum_45_1_2, cout_45_1_2;

full_adder fa_45_1_2(sum_45_1_2, cout_45_1_2, cout_44_3_1, cout_44_4_1, sum_45_0_1);

wire sum_45_2_2, cout_45_2_2;

full_adder fa_45_2_2(sum_45_2_2, cout_45_2_2, sum_45_1_1, sum_45_2_1, sum_45_3_1);

wire sum_46_0_2, cout_46_0_2;

full_adder fa_46_0_2(sum_46_0_2, cout_46_0_2, cout_45_0_1, cout_45_1_1, cout_45_2_1);

wire sum_46_1_2, cout_46_1_2;

full_adder fa_46_1_2(sum_46_1_2, cout_46_1_2, cout_45_3_1, sum_46_0_1, sum_46_1_1);

wire sum_46_2_2, cout_46_2_2;

half_adder ha_46_2_2(sum_46_2_2, cout_46_2_2, sum_46_2_1, sum_46_3_1);

wire sum_47_0_2, cout_47_0_2;

full_adder fa_47_0_2(sum_47_0_2, cout_47_0_2, cout_46_0_1, cout_46_1_1, cout_46_2_1);

wire sum_47_1_2, cout_47_1_2;

full_adder fa_47_1_2(sum_47_1_2, cout_47_1_2, cout_46_3_1, sum_47_0_1, sum_47_1_1);

wire sum_47_2_2, cout_47_2_2;

half_adder ha_47_2_2(sum_47_2_2, cout_47_2_2, sum_47_2_1, sum_47_3_1);

wire sum_48_0_2, cout_48_0_2;

full_adder fa_48_0_2(sum_48_0_2, cout_48_0_2, sum_48_4_0, cout_47_0_1, cout_47_1_1);

wire sum_48_1_2, cout_48_1_2;

full_adder fa_48_1_2(sum_48_1_2, cout_48_1_2, cout_47_2_1, cout_47_3_1, sum_48_0_1);

wire sum_48_2_2, cout_48_2_2;

half_adder ha_48_2_2(sum_48_2_2, cout_48_2_2, sum_48_1_1, sum_48_2_1);

wire sum_49_0_2, cout_49_0_2;

full_adder fa_49_0_2(sum_49_0_2, cout_49_0_2, sum_49_4_0, cout_48_0_1, cout_48_1_1);

wire sum_49_1_2, cout_49_1_2;

full_adder fa_49_1_2(sum_49_1_2, cout_49_1_2, cout_48_2_1, sum_49_0_1, sum_49_1_1);

wire sum_50_0_2, cout_50_0_2;

full_adder fa_50_0_2(sum_50_0_2, cout_50_0_2, sum_50_3_0, cout_49_0_1, cout_49_1_1);

wire sum_50_1_2, cout_50_1_2;

full_adder fa_50_1_2(sum_50_1_2, cout_50_1_2, cout_49_2_1, sum_50_0_1, sum_50_1_1);

wire sum_51_0_2, cout_51_0_2;

full_adder fa_51_0_2(sum_51_0_2, cout_51_0_2, cout_50_0_1, cout_50_1_1, cout_50_2_1);

wire sum_51_1_2, cout_51_1_2;

full_adder fa_51_1_2(sum_51_1_2, cout_51_1_2, sum_51_0_1, sum_51_1_1, sum_51_2_1);

wire sum_52_0_2, cout_52_0_2;

full_adder fa_52_0_2(sum_52_0_2, cout_52_0_2, cout_51_0_1, cout_51_1_1, cout_51_2_1);

wire sum_52_1_2, cout_52_1_2;

full_adder fa_52_1_2(sum_52_1_2, cout_52_1_2, sum_52_0_1, sum_52_1_1, sum_52_2_1);

wire sum_53_0_2, cout_53_0_2;

full_adder fa_53_0_2(sum_53_0_2, cout_53_0_2, cout_52_0_1, cout_52_1_1, cout_52_2_1);

wire sum_53_1_2, cout_53_1_2;

full_adder fa_53_1_2(sum_53_1_2, cout_53_1_2, sum_53_0_1, sum_53_1_1, sum_53_2_1);

wire sum_54_0_2, cout_54_0_2;

full_adder fa_54_0_2(sum_54_0_2, cout_54_0_2, cout_53_0_1, cout_53_1_1, cout_53_2_1);

wire sum_54_1_2, cout_54_1_2;

half_adder ha_54_1_2(sum_54_1_2, cout_54_1_2, sum_54_0_1, sum_54_1_1);

wire sum_55_0_2, cout_55_0_2;

full_adder fa_55_0_2(sum_55_0_2, cout_55_0_2, cout_54_0_1, cout_54_1_1, sum_55_0_1);

wire sum_56_0_2, cout_56_0_2;

full_adder fa_56_0_2(sum_56_0_2, cout_56_0_2, cout_55_0_1, cout_55_1_1, sum_56_0_1);

wire sum_57_0_2, cout_57_0_2;

full_adder fa_57_0_2(sum_57_0_2, cout_57_0_2, sum_57_1_0, cout_56_0_1, cout_56_1_1);

wire sum_58_0_2, cout_58_0_2;

full_adder fa_58_0_2(sum_58_0_2, cout_58_0_2, sum_58_1_0, cout_57_0_1, sum_58_0_1);

wire sum_59_0_2, cout_59_0_2;

full_adder fa_59_0_2(sum_59_0_2, cout_59_0_2, sum_59_0_0, cout_58_0_1, sum_59_0_1);

wire sum_60_0_2, cout_60_0_2;

full_adder fa_60_0_2(sum_60_0_2, cout_60_0_2, cout_59_0_0, sum_60_0_0, cout_59_0_1);

wire sum_61_0_2, cout_61_0_2;

full_adder fa_61_0_2(sum_61_0_2, cout_61_0_2, A31B30, A30B31, cout_60_0_0);

wire sum_7_0_3, cout_7_0_3;

half_adder ha_7_0_3(sum_7_0_3, cout_7_0_3, sum_7_1_1, cout_6_0_2);

wire sum_8_0_3, cout_8_0_3;

full_adder fa_8_0_3(sum_8_0_3, cout_8_0_3, sum_8_1_1, cout_7_0_2, sum_8_0_2);

wire sum_9_0_3, cout_9_0_3;

full_adder fa_9_0_3(sum_9_0_3, cout_9_0_3, cout_8_0_2, sum_9_0_2, sum_9_1_2);

wire sum_10_0_3, cout_10_0_3;

full_adder fa_10_0_3(sum_10_0_3, cout_10_0_3, cout_9_0_2, cout_9_1_2, sum_10_0_2);

wire sum_11_0_3, cout_11_0_3;

full_adder fa_11_0_3(sum_11_0_3, cout_11_0_3, cout_10_0_2, cout_10_1_2, sum_11_0_2);

wire sum_12_0_3, cout_12_0_3;

full_adder fa_12_0_3(sum_12_0_3, cout_12_0_3, cout_11_0_2, cout_11_1_2, sum_12_0_2);

wire sum_13_0_3, cout_13_0_3;

full_adder fa_13_0_3(sum_13_0_3, cout_13_0_3, cout_12_0_2, cout_12_1_2, sum_13_0_2);

wire sum_14_0_3, cout_14_0_3;

full_adder fa_14_0_3(sum_14_0_3, cout_14_0_3, sum_14_2_1, cout_13_0_2, cout_13_1_2);

wire sum_14_1_3, cout_14_1_3;

half_adder ha_14_1_3(sum_14_1_3, cout_14_1_3, sum_14_0_2, sum_14_1_2);

wire sum_15_0_3, cout_15_0_3;

full_adder fa_15_0_3(sum_15_0_3, cout_15_0_3, sum_15_3_1, cout_14_0_2, cout_14_1_2);

wire sum_15_1_3, cout_15_1_3;

half_adder ha_15_1_3(sum_15_1_3, cout_15_1_3, sum_15_0_2, sum_15_1_2);

wire sum_16_0_3, cout_16_0_3;

full_adder fa_16_0_3(sum_16_0_3, cout_16_0_3, cout_15_0_2, cout_15_1_2, sum_16_0_2);

wire sum_16_1_3, cout_16_1_3;

half_adder ha_16_1_3(sum_16_1_3, cout_16_1_3, sum_16_1_2, sum_16_2_2);

wire sum_17_0_3, cout_17_0_3;

full_adder fa_17_0_3(sum_17_0_3, cout_17_0_3, cout_16_0_2, cout_16_1_2, cout_16_2_2);

wire sum_17_1_3, cout_17_1_3;

full_adder fa_17_1_3(sum_17_1_3, cout_17_1_3, sum_17_0_2, sum_17_1_2, sum_17_2_2);

wire sum_18_0_3, cout_18_0_3;

full_adder fa_18_0_3(sum_18_0_3, cout_18_0_3, cout_17_0_2, cout_17_1_2, cout_17_2_2);

wire sum_18_1_3, cout_18_1_3;

full_adder fa_18_1_3(sum_18_1_3, cout_18_1_3, sum_18_0_2, sum_18_1_2, sum_18_2_2);

wire sum_19_0_3, cout_19_0_3;

full_adder fa_19_0_3(sum_19_0_3, cout_19_0_3, cout_18_0_2, cout_18_1_2, cout_18_2_2);

wire sum_19_1_3, cout_19_1_3;

full_adder fa_19_1_3(sum_19_1_3, cout_19_1_3, sum_19_0_2, sum_19_1_2, sum_19_2_2);

wire sum_20_0_3, cout_20_0_3;

full_adder fa_20_0_3(sum_20_0_3, cout_20_0_3, cout_19_0_2, cout_19_1_2, cout_19_2_2);

wire sum_20_1_3, cout_20_1_3;

full_adder fa_20_1_3(sum_20_1_3, cout_20_1_3, sum_20_0_2, sum_20_1_2, sum_20_2_2);

wire sum_21_0_3, cout_21_0_3;

full_adder fa_21_0_3(sum_21_0_3, cout_21_0_3, sum_21_4_1, cout_20_0_2, cout_20_1_2);

wire sum_21_1_3, cout_21_1_3;

full_adder fa_21_1_3(sum_21_1_3, cout_21_1_3, cout_20_2_2, sum_21_0_2, sum_21_1_2);

wire sum_22_0_3, cout_22_0_3;

full_adder fa_22_0_3(sum_22_0_3, cout_22_0_3, sum_22_4_1, cout_21_0_2, cout_21_1_2);

wire sum_22_1_3, cout_22_1_3;

full_adder fa_22_1_3(sum_22_1_3, cout_22_1_3, cout_21_2_2, sum_22_0_2, sum_22_1_2);

wire sum_23_0_3, cout_23_0_3;

full_adder fa_23_0_3(sum_23_0_3, cout_23_0_3, cout_22_0_2, cout_22_1_2, cout_22_2_2);

wire sum_23_1_3, cout_23_1_3;

full_adder fa_23_1_3(sum_23_1_3, cout_23_1_3, sum_23_0_2, sum_23_1_2, sum_23_2_2);

wire sum_24_0_3, cout_24_0_3;

full_adder fa_24_0_3(sum_24_0_3, cout_24_0_3, cout_23_0_2, cout_23_1_2, cout_23_2_2);

wire sum_24_1_3, cout_24_1_3;

full_adder fa_24_1_3(sum_24_1_3, cout_24_1_3, cout_23_3_2, sum_24_0_2, sum_24_1_2);

wire sum_24_2_3, cout_24_2_3;

half_adder ha_24_2_3(sum_24_2_3, cout_24_2_3, sum_24_2_2, sum_24_3_2);

wire sum_25_0_3, cout_25_0_3;

full_adder fa_25_0_3(sum_25_0_3, cout_25_0_3, cout_24_0_2, cout_24_1_2, cout_24_2_2);

wire sum_25_1_3, cout_25_1_3;

full_adder fa_25_1_3(sum_25_1_3, cout_25_1_3, cout_24_3_2, sum_25_0_2, sum_25_1_2);

wire sum_25_2_3, cout_25_2_3;

half_adder ha_25_2_3(sum_25_2_3, cout_25_2_3, sum_25_2_2, sum_25_3_2);

wire sum_26_0_3, cout_26_0_3;

full_adder fa_26_0_3(sum_26_0_3, cout_26_0_3, cout_25_0_2, cout_25_1_2, cout_25_2_2);

wire sum_26_1_3, cout_26_1_3;

full_adder fa_26_1_3(sum_26_1_3, cout_26_1_3, cout_25_3_2, sum_26_0_2, sum_26_1_2);

wire sum_26_2_3, cout_26_2_3;

half_adder ha_26_2_3(sum_26_2_3, cout_26_2_3, sum_26_2_2, sum_26_3_2);

wire sum_27_0_3, cout_27_0_3;

full_adder fa_27_0_3(sum_27_0_3, cout_27_0_3, sum_27_5_1, cout_26_0_2, cout_26_1_2);

wire sum_27_1_3, cout_27_1_3;

full_adder fa_27_1_3(sum_27_1_3, cout_27_1_3, cout_26_2_2, cout_26_3_2, sum_27_0_2);

wire sum_27_2_3, cout_27_2_3;

full_adder fa_27_2_3(sum_27_2_3, cout_27_2_3, sum_27_1_2, sum_27_2_2, sum_27_3_2);

wire sum_28_0_3, cout_28_0_3;

full_adder fa_28_0_3(sum_28_0_3, cout_28_0_3, sum_28_5_1, cout_27_0_2, cout_27_1_2);

wire sum_28_1_3, cout_28_1_3;

full_adder fa_28_1_3(sum_28_1_3, cout_28_1_3, cout_27_2_2, cout_27_3_2, sum_28_0_2);

wire sum_28_2_3, cout_28_2_3;

full_adder fa_28_2_3(sum_28_2_3, cout_28_2_3, sum_28_1_2, sum_28_2_2, sum_28_3_2);

wire sum_29_0_3, cout_29_0_3;

full_adder fa_29_0_3(sum_29_0_3, cout_29_0_3, sum_29_6_1, cout_28_0_2, cout_28_1_2);

wire sum_29_1_3, cout_29_1_3;

full_adder fa_29_1_3(sum_29_1_3, cout_29_1_3, cout_28_2_2, cout_28_3_2, sum_29_0_2);

wire sum_29_2_3, cout_29_2_3;

full_adder fa_29_2_3(sum_29_2_3, cout_29_2_3, sum_29_1_2, sum_29_2_2, sum_29_3_2);

wire sum_30_0_3, cout_30_0_3;

full_adder fa_30_0_3(sum_30_0_3, cout_30_0_3, cout_29_0_2, cout_29_1_2, cout_29_2_2);

wire sum_30_1_3, cout_30_1_3;

full_adder fa_30_1_3(sum_30_1_3, cout_30_1_3, cout_29_3_2, sum_30_0_2, sum_30_1_2);

wire sum_30_2_3, cout_30_2_3;

full_adder fa_30_2_3(sum_30_2_3, cout_30_2_3, sum_30_2_2, sum_30_3_2, sum_30_4_2);

wire sum_31_0_3, cout_31_0_3;

full_adder fa_31_0_3(sum_31_0_3, cout_31_0_3, cout_30_0_2, cout_30_1_2, cout_30_2_2);

wire sum_31_1_3, cout_31_1_3;

full_adder fa_31_1_3(sum_31_1_3, cout_31_1_3, cout_30_3_2, cout_30_4_2, sum_31_0_2);

wire sum_31_2_3, cout_31_2_3;

full_adder fa_31_2_3(sum_31_2_3, cout_31_2_3, sum_31_1_2, sum_31_2_2, sum_31_3_2);

wire sum_32_0_3, cout_32_0_3;

full_adder fa_32_0_3(sum_32_0_3, cout_32_0_3, cout_31_0_2, cout_31_1_2, cout_31_2_2);

wire sum_32_1_3, cout_32_1_3;

full_adder fa_32_1_3(sum_32_1_3, cout_32_1_3, cout_31_3_2, cout_31_4_2, sum_32_0_2);

wire sum_32_2_3, cout_32_2_3;

full_adder fa_32_2_3(sum_32_2_3, cout_32_2_3, sum_32_1_2, sum_32_2_2, sum_32_3_2);

wire sum_33_0_3, cout_33_0_3;

full_adder fa_33_0_3(sum_33_0_3, cout_33_0_3, cout_32_0_2, cout_32_1_2, cout_32_2_2);

wire sum_33_1_3, cout_33_1_3;

full_adder fa_33_1_3(sum_33_1_3, cout_33_1_3, cout_32_3_2, cout_32_4_2, sum_33_0_2);

wire sum_33_2_3, cout_33_2_3;

full_adder fa_33_2_3(sum_33_2_3, cout_33_2_3, sum_33_1_2, sum_33_2_2, sum_33_3_2);

wire sum_34_0_3, cout_34_0_3;

full_adder fa_34_0_3(sum_34_0_3, cout_34_0_3, cout_33_0_2, cout_33_1_2, cout_33_2_2);

wire sum_34_1_3, cout_34_1_3;

full_adder fa_34_1_3(sum_34_1_3, cout_34_1_3, cout_33_3_2, cout_33_4_2, sum_34_0_2);

wire sum_34_2_3, cout_34_2_3;

full_adder fa_34_2_3(sum_34_2_3, cout_34_2_3, sum_34_1_2, sum_34_2_2, sum_34_3_2);

wire sum_35_0_3, cout_35_0_3;

full_adder fa_35_0_3(sum_35_0_3, cout_35_0_3, cout_34_0_2, cout_34_1_2, cout_34_2_2);

wire sum_35_1_3, cout_35_1_3;

full_adder fa_35_1_3(sum_35_1_3, cout_35_1_3, cout_34_3_2, cout_34_4_2, sum_35_0_2);

wire sum_35_2_3, cout_35_2_3;

full_adder fa_35_2_3(sum_35_2_3, cout_35_2_3, sum_35_1_2, sum_35_2_2, sum_35_3_2);

wire sum_36_0_3, cout_36_0_3;

full_adder fa_36_0_3(sum_36_0_3, cout_36_0_3, sum_36_5_1, cout_35_0_2, cout_35_1_2);

wire sum_36_1_3, cout_36_1_3;

full_adder fa_36_1_3(sum_36_1_3, cout_36_1_3, cout_35_2_2, cout_35_3_2, cout_35_4_2);

wire sum_36_2_3, cout_36_2_3;

full_adder fa_36_2_3(sum_36_2_3, cout_36_2_3, sum_36_0_2, sum_36_1_2, sum_36_2_2);

wire sum_37_0_3, cout_37_0_3;

full_adder fa_37_0_3(sum_37_0_3, cout_37_0_3, cout_36_0_2, cout_36_1_2, cout_36_2_2);

wire sum_37_1_3, cout_37_1_3;

full_adder fa_37_1_3(sum_37_1_3, cout_37_1_3, cout_36_3_2, sum_37_0_2, sum_37_1_2);

wire sum_37_2_3, cout_37_2_3;

half_adder ha_37_2_3(sum_37_2_3, cout_37_2_3, sum_37_2_2, sum_37_3_2);

wire sum_38_0_3, cout_38_0_3;

full_adder fa_38_0_3(sum_38_0_3, cout_38_0_3, cout_37_0_2, cout_37_1_2, cout_37_2_2);

wire sum_38_1_3, cout_38_1_3;

full_adder fa_38_1_3(sum_38_1_3, cout_38_1_3, cout_37_3_2, sum_38_0_2, sum_38_1_2);

wire sum_38_2_3, cout_38_2_3;

half_adder ha_38_2_3(sum_38_2_3, cout_38_2_3, sum_38_2_2, sum_38_3_2);

wire sum_39_0_3, cout_39_0_3;

full_adder fa_39_0_3(sum_39_0_3, cout_39_0_3, cout_38_0_2, cout_38_1_2, cout_38_2_2);

wire sum_39_1_3, cout_39_1_3;

full_adder fa_39_1_3(sum_39_1_3, cout_39_1_3, cout_38_3_2, sum_39_0_2, sum_39_1_2);

wire sum_39_2_3, cout_39_2_3;

half_adder ha_39_2_3(sum_39_2_3, cout_39_2_3, sum_39_2_2, sum_39_3_2);

wire sum_40_0_3, cout_40_0_3;

full_adder fa_40_0_3(sum_40_0_3, cout_40_0_3, cout_39_0_2, cout_39_1_2, cout_39_2_2);

wire sum_40_1_3, cout_40_1_3;

full_adder fa_40_1_3(sum_40_1_3, cout_40_1_3, cout_39_3_2, sum_40_0_2, sum_40_1_2);

wire sum_40_2_3, cout_40_2_3;

half_adder ha_40_2_3(sum_40_2_3, cout_40_2_3, sum_40_2_2, sum_40_3_2);

wire sum_41_0_3, cout_41_0_3;

full_adder fa_41_0_3(sum_41_0_3, cout_41_0_3, cout_40_0_2, cout_40_1_2, cout_40_2_2);

wire sum_41_1_3, cout_41_1_3;

full_adder fa_41_1_3(sum_41_1_3, cout_41_1_3, cout_40_3_2, sum_41_0_2, sum_41_1_2);

wire sum_41_2_3, cout_41_2_3;

half_adder ha_41_2_3(sum_41_2_3, cout_41_2_3, sum_41_2_2, sum_41_3_2);

wire sum_42_0_3, cout_42_0_3;

full_adder fa_42_0_3(sum_42_0_3, cout_42_0_3, sum_42_4_1, cout_41_0_2, cout_41_1_2);

wire sum_42_1_3, cout_42_1_3;

full_adder fa_42_1_3(sum_42_1_3, cout_42_1_3, cout_41_2_2, cout_41_3_2, sum_42_0_2);

wire sum_42_2_3, cout_42_2_3;

half_adder ha_42_2_3(sum_42_2_3, cout_42_2_3, sum_42_1_2, sum_42_2_2);

wire sum_43_0_3, cout_43_0_3;

full_adder fa_43_0_3(sum_43_0_3, cout_43_0_3, sum_43_4_1, cout_42_0_2, cout_42_1_2);

wire sum_43_1_3, cout_43_1_3;

full_adder fa_43_1_3(sum_43_1_3, cout_43_1_3, cout_42_2_2, sum_43_0_2, sum_43_1_2);

wire sum_44_0_3, cout_44_0_3;

full_adder fa_44_0_3(sum_44_0_3, cout_44_0_3, sum_44_4_1, cout_43_0_2, cout_43_1_2);

wire sum_44_1_3, cout_44_1_3;

full_adder fa_44_1_3(sum_44_1_3, cout_44_1_3, cout_43_2_2, sum_44_0_2, sum_44_1_2);

wire sum_45_0_3, cout_45_0_3;

full_adder fa_45_0_3(sum_45_0_3, cout_45_0_3, cout_44_0_2, cout_44_1_2, cout_44_2_2);

wire sum_45_1_3, cout_45_1_3;

full_adder fa_45_1_3(sum_45_1_3, cout_45_1_3, sum_45_0_2, sum_45_1_2, sum_45_2_2);

wire sum_46_0_3, cout_46_0_3;

full_adder fa_46_0_3(sum_46_0_3, cout_46_0_3, cout_45_0_2, cout_45_1_2, cout_45_2_2);

wire sum_46_1_3, cout_46_1_3;

full_adder fa_46_1_3(sum_46_1_3, cout_46_1_3, sum_46_0_2, sum_46_1_2, sum_46_2_2);

wire sum_47_0_3, cout_47_0_3;

full_adder fa_47_0_3(sum_47_0_3, cout_47_0_3, cout_46_0_2, cout_46_1_2, cout_46_2_2);

wire sum_47_1_3, cout_47_1_3;

full_adder fa_47_1_3(sum_47_1_3, cout_47_1_3, sum_47_0_2, sum_47_1_2, sum_47_2_2);

wire sum_48_0_3, cout_48_0_3;

full_adder fa_48_0_3(sum_48_0_3, cout_48_0_3, cout_47_0_2, cout_47_1_2, cout_47_2_2);

wire sum_48_1_3, cout_48_1_3;

full_adder fa_48_1_3(sum_48_1_3, cout_48_1_3, sum_48_0_2, sum_48_1_2, sum_48_2_2);

wire sum_49_0_3, cout_49_0_3;

full_adder fa_49_0_3(sum_49_0_3, cout_49_0_3, sum_49_2_1, cout_48_0_2, cout_48_1_2);

wire sum_49_1_3, cout_49_1_3;

full_adder fa_49_1_3(sum_49_1_3, cout_49_1_3, cout_48_2_2, sum_49_0_2, sum_49_1_2);

wire sum_50_0_3, cout_50_0_3;

full_adder fa_50_0_3(sum_50_0_3, cout_50_0_3, sum_50_2_1, cout_49_0_2, cout_49_1_2);

wire sum_50_1_3, cout_50_1_3;

half_adder ha_50_1_3(sum_50_1_3, cout_50_1_3, sum_50_0_2, sum_50_1_2);

wire sum_51_0_3, cout_51_0_3;

full_adder fa_51_0_3(sum_51_0_3, cout_51_0_3, cout_50_0_2, cout_50_1_2, sum_51_0_2);

wire sum_52_0_3, cout_52_0_3;

full_adder fa_52_0_3(sum_52_0_3, cout_52_0_3, cout_51_0_2, cout_51_1_2, sum_52_0_2);

wire sum_53_0_3, cout_53_0_3;

full_adder fa_53_0_3(sum_53_0_3, cout_53_0_3, cout_52_0_2, cout_52_1_2, sum_53_0_2);

wire sum_54_0_3, cout_54_0_3;

full_adder fa_54_0_3(sum_54_0_3, cout_54_0_3, cout_53_0_2, cout_53_1_2, sum_54_0_2);

wire sum_55_0_3, cout_55_0_3;

full_adder fa_55_0_3(sum_55_0_3, cout_55_0_3, sum_55_1_1, cout_54_0_2, cout_54_1_2);

wire sum_56_0_3, cout_56_0_3;

full_adder fa_56_0_3(sum_56_0_3, cout_56_0_3, sum_56_1_1, cout_55_0_2, sum_56_0_2);

wire sum_57_0_3, cout_57_0_3;

full_adder fa_57_0_3(sum_57_0_3, cout_57_0_3, sum_57_0_1, cout_56_0_2, sum_57_0_2);

wire sum_10_0_4, cout_10_0_4;

half_adder ha_10_0_4(sum_10_0_4, cout_10_0_4, sum_10_1_2, cout_9_0_3);

wire sum_11_0_4, cout_11_0_4;

full_adder fa_11_0_4(sum_11_0_4, cout_11_0_4, sum_11_1_2, cout_10_0_3, sum_11_0_3);

wire sum_12_0_4, cout_12_0_4;

full_adder fa_12_0_4(sum_12_0_4, cout_12_0_4, sum_12_1_2, cout_11_0_3, sum_12_0_3);

wire sum_13_0_4, cout_13_0_4;

full_adder fa_13_0_4(sum_13_0_4, cout_13_0_4, sum_13_1_2, cout_12_0_3, sum_13_0_3);

wire sum_14_0_4, cout_14_0_4;

full_adder fa_14_0_4(sum_14_0_4, cout_14_0_4, cout_13_0_3, sum_14_0_3, sum_14_1_3);

wire sum_15_0_4, cout_15_0_4;

full_adder fa_15_0_4(sum_15_0_4, cout_15_0_4, cout_14_0_3, cout_14_1_3, sum_15_0_3);

wire sum_16_0_4, cout_16_0_4;

full_adder fa_16_0_4(sum_16_0_4, cout_16_0_4, cout_15_0_3, cout_15_1_3, sum_16_0_3);

wire sum_17_0_4, cout_17_0_4;

full_adder fa_17_0_4(sum_17_0_4, cout_17_0_4, cout_16_0_3, cout_16_1_3, sum_17_0_3);

wire sum_18_0_4, cout_18_0_4;

full_adder fa_18_0_4(sum_18_0_4, cout_18_0_4, cout_17_0_3, cout_17_1_3, sum_18_0_3);

wire sum_19_0_4, cout_19_0_4;

full_adder fa_19_0_4(sum_19_0_4, cout_19_0_4, cout_18_0_3, cout_18_1_3, sum_19_0_3);

wire sum_20_0_4, cout_20_0_4;

full_adder fa_20_0_4(sum_20_0_4, cout_20_0_4, cout_19_0_3, cout_19_1_3, sum_20_0_3);

wire sum_21_0_4, cout_21_0_4;

full_adder fa_21_0_4(sum_21_0_4, cout_21_0_4, sum_21_2_2, cout_20_0_3, cout_20_1_3);

wire sum_21_1_4, cout_21_1_4;

half_adder ha_21_1_4(sum_21_1_4, cout_21_1_4, sum_21_0_3, sum_21_1_3);

wire sum_22_0_4, cout_22_0_4;

full_adder fa_22_0_4(sum_22_0_4, cout_22_0_4, sum_22_2_2, cout_21_0_3, cout_21_1_3);

wire sum_22_1_4, cout_22_1_4;

half_adder ha_22_1_4(sum_22_1_4, cout_22_1_4, sum_22_0_3, sum_22_1_3);

wire sum_23_0_4, cout_23_0_4;

full_adder fa_23_0_4(sum_23_0_4, cout_23_0_4, sum_23_3_2, cout_22_0_3, cout_22_1_3);

wire sum_23_1_4, cout_23_1_4;

half_adder ha_23_1_4(sum_23_1_4, cout_23_1_4, sum_23_0_3, sum_23_1_3);

wire sum_24_0_4, cout_24_0_4;

full_adder fa_24_0_4(sum_24_0_4, cout_24_0_4, cout_23_0_3, cout_23_1_3, sum_24_0_3);

wire sum_24_1_4, cout_24_1_4;

half_adder ha_24_1_4(sum_24_1_4, cout_24_1_4, sum_24_1_3, sum_24_2_3);

wire sum_25_0_4, cout_25_0_4;

full_adder fa_25_0_4(sum_25_0_4, cout_25_0_4, cout_24_0_3, cout_24_1_3, cout_24_2_3);

wire sum_25_1_4, cout_25_1_4;

full_adder fa_25_1_4(sum_25_1_4, cout_25_1_4, sum_25_0_3, sum_25_1_3, sum_25_2_3);

wire sum_26_0_4, cout_26_0_4;

full_adder fa_26_0_4(sum_26_0_4, cout_26_0_4, cout_25_0_3, cout_25_1_3, cout_25_2_3);

wire sum_26_1_4, cout_26_1_4;

full_adder fa_26_1_4(sum_26_1_4, cout_26_1_4, sum_26_0_3, sum_26_1_3, sum_26_2_3);

wire sum_27_0_4, cout_27_0_4;

full_adder fa_27_0_4(sum_27_0_4, cout_27_0_4, cout_26_0_3, cout_26_1_3, cout_26_2_3);

wire sum_27_1_4, cout_27_1_4;

full_adder fa_27_1_4(sum_27_1_4, cout_27_1_4, sum_27_0_3, sum_27_1_3, sum_27_2_3);

wire sum_28_0_4, cout_28_0_4;

full_adder fa_28_0_4(sum_28_0_4, cout_28_0_4, cout_27_0_3, cout_27_1_3, cout_27_2_3);

wire sum_28_1_4, cout_28_1_4;

full_adder fa_28_1_4(sum_28_1_4, cout_28_1_4, sum_28_0_3, sum_28_1_3, sum_28_2_3);

wire sum_29_0_4, cout_29_0_4;

full_adder fa_29_0_4(sum_29_0_4, cout_29_0_4, cout_28_0_3, cout_28_1_3, cout_28_2_3);

wire sum_29_1_4, cout_29_1_4;

full_adder fa_29_1_4(sum_29_1_4, cout_29_1_4, sum_29_0_3, sum_29_1_3, sum_29_2_3);

wire sum_30_0_4, cout_30_0_4;

full_adder fa_30_0_4(sum_30_0_4, cout_30_0_4, cout_29_0_3, cout_29_1_3, cout_29_2_3);

wire sum_30_1_4, cout_30_1_4;

full_adder fa_30_1_4(sum_30_1_4, cout_30_1_4, sum_30_0_3, sum_30_1_3, sum_30_2_3);

wire sum_31_0_4, cout_31_0_4;

full_adder fa_31_0_4(sum_31_0_4, cout_31_0_4, sum_31_4_2, cout_30_0_3, cout_30_1_3);

wire sum_31_1_4, cout_31_1_4;

full_adder fa_31_1_4(sum_31_1_4, cout_31_1_4, cout_30_2_3, sum_31_0_3, sum_31_1_3);

wire sum_32_0_4, cout_32_0_4;

full_adder fa_32_0_4(sum_32_0_4, cout_32_0_4, sum_32_4_2, cout_31_0_3, cout_31_1_3);

wire sum_32_1_4, cout_32_1_4;

full_adder fa_32_1_4(sum_32_1_4, cout_32_1_4, cout_31_2_3, sum_32_0_3, sum_32_1_3);

wire sum_33_0_4, cout_33_0_4;

full_adder fa_33_0_4(sum_33_0_4, cout_33_0_4, sum_33_4_2, cout_32_0_3, cout_32_1_3);

wire sum_33_1_4, cout_33_1_4;

full_adder fa_33_1_4(sum_33_1_4, cout_33_1_4, cout_32_2_3, sum_33_0_3, sum_33_1_3);

wire sum_34_0_4, cout_34_0_4;

full_adder fa_34_0_4(sum_34_0_4, cout_34_0_4, sum_34_4_2, cout_33_0_3, cout_33_1_3);

wire sum_34_1_4, cout_34_1_4;

full_adder fa_34_1_4(sum_34_1_4, cout_34_1_4, cout_33_2_3, sum_34_0_3, sum_34_1_3);

wire sum_35_0_4, cout_35_0_4;

full_adder fa_35_0_4(sum_35_0_4, cout_35_0_4, sum_35_4_2, cout_34_0_3, cout_34_1_3);

wire sum_35_1_4, cout_35_1_4;

full_adder fa_35_1_4(sum_35_1_4, cout_35_1_4, cout_34_2_3, sum_35_0_3, sum_35_1_3);

wire sum_36_0_4, cout_36_0_4;

full_adder fa_36_0_4(sum_36_0_4, cout_36_0_4, sum_36_3_2, cout_35_0_3, cout_35_1_3);

wire sum_36_1_4, cout_36_1_4;

full_adder fa_36_1_4(sum_36_1_4, cout_36_1_4, cout_35_2_3, sum_36_0_3, sum_36_1_3);

wire sum_37_0_4, cout_37_0_4;

full_adder fa_37_0_4(sum_37_0_4, cout_37_0_4, cout_36_0_3, cout_36_1_3, cout_36_2_3);

wire sum_37_1_4, cout_37_1_4;

full_adder fa_37_1_4(sum_37_1_4, cout_37_1_4, sum_37_0_3, sum_37_1_3, sum_37_2_3);

wire sum_38_0_4, cout_38_0_4;

full_adder fa_38_0_4(sum_38_0_4, cout_38_0_4, cout_37_0_3, cout_37_1_3, cout_37_2_3);

wire sum_38_1_4, cout_38_1_4;

full_adder fa_38_1_4(sum_38_1_4, cout_38_1_4, sum_38_0_3, sum_38_1_3, sum_38_2_3);

wire sum_39_0_4, cout_39_0_4;

full_adder fa_39_0_4(sum_39_0_4, cout_39_0_4, cout_38_0_3, cout_38_1_3, cout_38_2_3);

wire sum_39_1_4, cout_39_1_4;

full_adder fa_39_1_4(sum_39_1_4, cout_39_1_4, sum_39_0_3, sum_39_1_3, sum_39_2_3);

wire sum_40_0_4, cout_40_0_4;

full_adder fa_40_0_4(sum_40_0_4, cout_40_0_4, cout_39_0_3, cout_39_1_3, cout_39_2_3);

wire sum_40_1_4, cout_40_1_4;

full_adder fa_40_1_4(sum_40_1_4, cout_40_1_4, sum_40_0_3, sum_40_1_3, sum_40_2_3);

wire sum_41_0_4, cout_41_0_4;

full_adder fa_41_0_4(sum_41_0_4, cout_41_0_4, cout_40_0_3, cout_40_1_3, cout_40_2_3);

wire sum_41_1_4, cout_41_1_4;

full_adder fa_41_1_4(sum_41_1_4, cout_41_1_4, sum_41_0_3, sum_41_1_3, sum_41_2_3);

wire sum_42_0_4, cout_42_0_4;

full_adder fa_42_0_4(sum_42_0_4, cout_42_0_4, cout_41_0_3, cout_41_1_3, cout_41_2_3);

wire sum_42_1_4, cout_42_1_4;

full_adder fa_42_1_4(sum_42_1_4, cout_42_1_4, sum_42_0_3, sum_42_1_3, sum_42_2_3);

wire sum_43_0_4, cout_43_0_4;

full_adder fa_43_0_4(sum_43_0_4, cout_43_0_4, sum_43_2_2, cout_42_0_3, cout_42_1_3);

wire sum_43_1_4, cout_43_1_4;

full_adder fa_43_1_4(sum_43_1_4, cout_43_1_4, cout_42_2_3, sum_43_0_3, sum_43_1_3);

wire sum_44_0_4, cout_44_0_4;

full_adder fa_44_0_4(sum_44_0_4, cout_44_0_4, sum_44_2_2, cout_43_0_3, cout_43_1_3);

wire sum_44_1_4, cout_44_1_4;

half_adder ha_44_1_4(sum_44_1_4, cout_44_1_4, sum_44_0_3, sum_44_1_3);

wire sum_45_0_4, cout_45_0_4;

full_adder fa_45_0_4(sum_45_0_4, cout_45_0_4, cout_44_0_3, cout_44_1_3, sum_45_0_3);

wire sum_46_0_4, cout_46_0_4;

full_adder fa_46_0_4(sum_46_0_4, cout_46_0_4, cout_45_0_3, cout_45_1_3, sum_46_0_3);

wire sum_47_0_4, cout_47_0_4;

full_adder fa_47_0_4(sum_47_0_4, cout_47_0_4, cout_46_0_3, cout_46_1_3, sum_47_0_3);

wire sum_48_0_4, cout_48_0_4;

full_adder fa_48_0_4(sum_48_0_4, cout_48_0_4, cout_47_0_3, cout_47_1_3, sum_48_0_3);

wire sum_49_0_4, cout_49_0_4;

full_adder fa_49_0_4(sum_49_0_4, cout_49_0_4, cout_48_0_3, cout_48_1_3, sum_49_0_3);

wire sum_50_0_4, cout_50_0_4;

full_adder fa_50_0_4(sum_50_0_4, cout_50_0_4, cout_49_0_3, cout_49_1_3, sum_50_0_3);

wire sum_51_0_4, cout_51_0_4;

full_adder fa_51_0_4(sum_51_0_4, cout_51_0_4, sum_51_1_2, cout_50_0_3, cout_50_1_3);

wire sum_52_0_4, cout_52_0_4;

full_adder fa_52_0_4(sum_52_0_4, cout_52_0_4, sum_52_1_2, cout_51_0_3, sum_52_0_3);

wire sum_53_0_4, cout_53_0_4;

full_adder fa_53_0_4(sum_53_0_4, cout_53_0_4, sum_53_1_2, cout_52_0_3, sum_53_0_3);

wire sum_54_0_4, cout_54_0_4;

full_adder fa_54_0_4(sum_54_0_4, cout_54_0_4, sum_54_1_2, cout_53_0_3, sum_54_0_3);

wire sum_55_0_4, cout_55_0_4;

full_adder fa_55_0_4(sum_55_0_4, cout_55_0_4, sum_55_0_2, cout_54_0_3, sum_55_0_3);

wire sum_56_0_4, cout_56_0_4;

half_adder ha_56_0_4(sum_56_0_4, cout_56_0_4, cout_55_0_3, sum_56_0_3);

wire sum_57_0_4, cout_57_0_4;

half_adder ha_57_0_4(sum_57_0_4, cout_57_0_4, cout_56_0_3, sum_57_0_3);

wire sum_58_0_4, cout_58_0_4;

full_adder fa_58_0_4(sum_58_0_4, cout_58_0_4, cout_57_0_2, sum_58_0_2, cout_57_0_3);

wire sum_15_0_5, cout_15_0_5;

half_adder ha_15_0_5(sum_15_0_5, cout_15_0_5, sum_15_1_3, cout_14_0_4);

wire sum_16_0_5, cout_16_0_5;

full_adder fa_16_0_5(sum_16_0_5, cout_16_0_5, sum_16_1_3, cout_15_0_4, sum_16_0_4);

wire sum_17_0_5, cout_17_0_5;

full_adder fa_17_0_5(sum_17_0_5, cout_17_0_5, sum_17_1_3, cout_16_0_4, sum_17_0_4);

wire sum_18_0_5, cout_18_0_5;

full_adder fa_18_0_5(sum_18_0_5, cout_18_0_5, sum_18_1_3, cout_17_0_4, sum_18_0_4);

wire sum_19_0_5, cout_19_0_5;

full_adder fa_19_0_5(sum_19_0_5, cout_19_0_5, sum_19_1_3, cout_18_0_4, sum_19_0_4);

wire sum_20_0_5, cout_20_0_5;

full_adder fa_20_0_5(sum_20_0_5, cout_20_0_5, sum_20_1_3, cout_19_0_4, sum_20_0_4);

wire sum_21_0_5, cout_21_0_5;

full_adder fa_21_0_5(sum_21_0_5, cout_21_0_5, cout_20_0_4, sum_21_0_4, sum_21_1_4);

wire sum_22_0_5, cout_22_0_5;

full_adder fa_22_0_5(sum_22_0_5, cout_22_0_5, cout_21_0_4, cout_21_1_4, sum_22_0_4);

wire sum_23_0_5, cout_23_0_5;

full_adder fa_23_0_5(sum_23_0_5, cout_23_0_5, cout_22_0_4, cout_22_1_4, sum_23_0_4);

wire sum_24_0_5, cout_24_0_5;

full_adder fa_24_0_5(sum_24_0_5, cout_24_0_5, cout_23_0_4, cout_23_1_4, sum_24_0_4);

wire sum_25_0_5, cout_25_0_5;

full_adder fa_25_0_5(sum_25_0_5, cout_25_0_5, cout_24_0_4, cout_24_1_4, sum_25_0_4);

wire sum_26_0_5, cout_26_0_5;

full_adder fa_26_0_5(sum_26_0_5, cout_26_0_5, cout_25_0_4, cout_25_1_4, sum_26_0_4);

wire sum_27_0_5, cout_27_0_5;

full_adder fa_27_0_5(sum_27_0_5, cout_27_0_5, cout_26_0_4, cout_26_1_4, sum_27_0_4);

wire sum_28_0_5, cout_28_0_5;

full_adder fa_28_0_5(sum_28_0_5, cout_28_0_5, cout_27_0_4, cout_27_1_4, sum_28_0_4);

wire sum_29_0_5, cout_29_0_5;

full_adder fa_29_0_5(sum_29_0_5, cout_29_0_5, cout_28_0_4, cout_28_1_4, sum_29_0_4);

wire sum_30_0_5, cout_30_0_5;

full_adder fa_30_0_5(sum_30_0_5, cout_30_0_5, cout_29_0_4, cout_29_1_4, sum_30_0_4);

wire sum_31_0_5, cout_31_0_5;

full_adder fa_31_0_5(sum_31_0_5, cout_31_0_5, sum_31_2_3, cout_30_0_4, cout_30_1_4);

wire sum_31_1_5, cout_31_1_5;

half_adder ha_31_1_5(sum_31_1_5, cout_31_1_5, sum_31_0_4, sum_31_1_4);

wire sum_32_0_5, cout_32_0_5;

full_adder fa_32_0_5(sum_32_0_5, cout_32_0_5, sum_32_2_3, cout_31_0_4, cout_31_1_4);

wire sum_32_1_5, cout_32_1_5;

half_adder ha_32_1_5(sum_32_1_5, cout_32_1_5, sum_32_0_4, sum_32_1_4);

wire sum_33_0_5, cout_33_0_5;

full_adder fa_33_0_5(sum_33_0_5, cout_33_0_5, sum_33_2_3, cout_32_0_4, cout_32_1_4);

wire sum_33_1_5, cout_33_1_5;

half_adder ha_33_1_5(sum_33_1_5, cout_33_1_5, sum_33_0_4, sum_33_1_4);

wire sum_34_0_5, cout_34_0_5;

full_adder fa_34_0_5(sum_34_0_5, cout_34_0_5, sum_34_2_3, cout_33_0_4, cout_33_1_4);

wire sum_34_1_5, cout_34_1_5;

half_adder ha_34_1_5(sum_34_1_5, cout_34_1_5, sum_34_0_4, sum_34_1_4);

wire sum_35_0_5, cout_35_0_5;

full_adder fa_35_0_5(sum_35_0_5, cout_35_0_5, sum_35_2_3, cout_34_0_4, cout_34_1_4);

wire sum_35_1_5, cout_35_1_5;

half_adder ha_35_1_5(sum_35_1_5, cout_35_1_5, sum_35_0_4, sum_35_1_4);

wire sum_36_0_5, cout_36_0_5;

full_adder fa_36_0_5(sum_36_0_5, cout_36_0_5, sum_36_2_3, cout_35_0_4, cout_35_1_4);

wire sum_36_1_5, cout_36_1_5;

half_adder ha_36_1_5(sum_36_1_5, cout_36_1_5, sum_36_0_4, sum_36_1_4);

wire sum_37_0_5, cout_37_0_5;

full_adder fa_37_0_5(sum_37_0_5, cout_37_0_5, cout_36_0_4, cout_36_1_4, sum_37_0_4);

wire sum_38_0_5, cout_38_0_5;

full_adder fa_38_0_5(sum_38_0_5, cout_38_0_5, cout_37_0_4, cout_37_1_4, sum_38_0_4);

wire sum_39_0_5, cout_39_0_5;

full_adder fa_39_0_5(sum_39_0_5, cout_39_0_5, cout_38_0_4, cout_38_1_4, sum_39_0_4);

wire sum_40_0_5, cout_40_0_5;

full_adder fa_40_0_5(sum_40_0_5, cout_40_0_5, cout_39_0_4, cout_39_1_4, sum_40_0_4);

wire sum_41_0_5, cout_41_0_5;

full_adder fa_41_0_5(sum_41_0_5, cout_41_0_5, cout_40_0_4, cout_40_1_4, sum_41_0_4);

wire sum_42_0_5, cout_42_0_5;

full_adder fa_42_0_5(sum_42_0_5, cout_42_0_5, cout_41_0_4, cout_41_1_4, sum_42_0_4);

wire sum_43_0_5, cout_43_0_5;

full_adder fa_43_0_5(sum_43_0_5, cout_43_0_5, cout_42_0_4, cout_42_1_4, sum_43_0_4);

wire sum_44_0_5, cout_44_0_5;

full_adder fa_44_0_5(sum_44_0_5, cout_44_0_5, cout_43_0_4, cout_43_1_4, sum_44_0_4);

wire sum_45_0_5, cout_45_0_5;

full_adder fa_45_0_5(sum_45_0_5, cout_45_0_5, sum_45_1_3, cout_44_0_4, cout_44_1_4);

wire sum_46_0_5, cout_46_0_5;

full_adder fa_46_0_5(sum_46_0_5, cout_46_0_5, sum_46_1_3, cout_45_0_4, sum_46_0_4);

wire sum_47_0_5, cout_47_0_5;

full_adder fa_47_0_5(sum_47_0_5, cout_47_0_5, sum_47_1_3, cout_46_0_4, sum_47_0_4);

wire sum_48_0_5, cout_48_0_5;

full_adder fa_48_0_5(sum_48_0_5, cout_48_0_5, sum_48_1_3, cout_47_0_4, sum_48_0_4);

wire sum_49_0_5, cout_49_0_5;

full_adder fa_49_0_5(sum_49_0_5, cout_49_0_5, sum_49_1_3, cout_48_0_4, sum_49_0_4);

wire sum_50_0_5, cout_50_0_5;

full_adder fa_50_0_5(sum_50_0_5, cout_50_0_5, sum_50_1_3, cout_49_0_4, sum_50_0_4);

wire sum_51_0_5, cout_51_0_5;

full_adder fa_51_0_5(sum_51_0_5, cout_51_0_5, sum_51_0_3, cout_50_0_4, sum_51_0_4);

wire sum_52_0_5, cout_52_0_5;

half_adder ha_52_0_5(sum_52_0_5, cout_52_0_5, cout_51_0_4, sum_52_0_4);

wire sum_53_0_5, cout_53_0_5;

half_adder ha_53_0_5(sum_53_0_5, cout_53_0_5, cout_52_0_4, sum_53_0_4);

wire sum_54_0_5, cout_54_0_5;

half_adder ha_54_0_5(sum_54_0_5, cout_54_0_5, cout_53_0_4, sum_54_0_4);

wire sum_55_0_5, cout_55_0_5;

half_adder ha_55_0_5(sum_55_0_5, cout_55_0_5, cout_54_0_4, sum_55_0_4);

wire sum_56_0_5, cout_56_0_5;

half_adder ha_56_0_5(sum_56_0_5, cout_56_0_5, cout_55_0_4, sum_56_0_4);

wire sum_57_0_5, cout_57_0_5;

half_adder ha_57_0_5(sum_57_0_5, cout_57_0_5, cout_56_0_4, sum_57_0_4);

wire sum_58_0_5, cout_58_0_5;

half_adder ha_58_0_5(sum_58_0_5, cout_58_0_5, cout_57_0_4, sum_58_0_4);

wire sum_59_0_5, cout_59_0_5;

full_adder fa_59_0_5(sum_59_0_5, cout_59_0_5, cout_58_0_2, sum_59_0_2, cout_58_0_4);

wire sum_22_0_6, cout_22_0_6;

half_adder ha_22_0_6(sum_22_0_6, cout_22_0_6, sum_22_1_4, cout_21_0_5);

wire sum_23_0_6, cout_23_0_6;

full_adder fa_23_0_6(sum_23_0_6, cout_23_0_6, sum_23_1_4, cout_22_0_5, sum_23_0_5);

wire sum_24_0_6, cout_24_0_6;

full_adder fa_24_0_6(sum_24_0_6, cout_24_0_6, sum_24_1_4, cout_23_0_5, sum_24_0_5);

wire sum_25_0_6, cout_25_0_6;

full_adder fa_25_0_6(sum_25_0_6, cout_25_0_6, sum_25_1_4, cout_24_0_5, sum_25_0_5);

wire sum_26_0_6, cout_26_0_6;

full_adder fa_26_0_6(sum_26_0_6, cout_26_0_6, sum_26_1_4, cout_25_0_5, sum_26_0_5);

wire sum_27_0_6, cout_27_0_6;

full_adder fa_27_0_6(sum_27_0_6, cout_27_0_6, sum_27_1_4, cout_26_0_5, sum_27_0_5);

wire sum_28_0_6, cout_28_0_6;

full_adder fa_28_0_6(sum_28_0_6, cout_28_0_6, sum_28_1_4, cout_27_0_5, sum_28_0_5);

wire sum_29_0_6, cout_29_0_6;

full_adder fa_29_0_6(sum_29_0_6, cout_29_0_6, sum_29_1_4, cout_28_0_5, sum_29_0_5);

wire sum_30_0_6, cout_30_0_6;

full_adder fa_30_0_6(sum_30_0_6, cout_30_0_6, sum_30_1_4, cout_29_0_5, sum_30_0_5);

wire sum_31_0_6, cout_31_0_6;

full_adder fa_31_0_6(sum_31_0_6, cout_31_0_6, cout_30_0_5, sum_31_0_5, sum_31_1_5);

wire sum_32_0_6, cout_32_0_6;

full_adder fa_32_0_6(sum_32_0_6, cout_32_0_6, cout_31_0_5, cout_31_1_5, sum_32_0_5);

wire sum_33_0_6, cout_33_0_6;

full_adder fa_33_0_6(sum_33_0_6, cout_33_0_6, cout_32_0_5, cout_32_1_5, sum_33_0_5);

wire sum_34_0_6, cout_34_0_6;

full_adder fa_34_0_6(sum_34_0_6, cout_34_0_6, cout_33_0_5, cout_33_1_5, sum_34_0_5);

wire sum_35_0_6, cout_35_0_6;

full_adder fa_35_0_6(sum_35_0_6, cout_35_0_6, cout_34_0_5, cout_34_1_5, sum_35_0_5);

wire sum_36_0_6, cout_36_0_6;

full_adder fa_36_0_6(sum_36_0_6, cout_36_0_6, cout_35_0_5, cout_35_1_5, sum_36_0_5);

wire sum_37_0_6, cout_37_0_6;

full_adder fa_37_0_6(sum_37_0_6, cout_37_0_6, sum_37_1_4, cout_36_0_5, cout_36_1_5);

wire sum_38_0_6, cout_38_0_6;

full_adder fa_38_0_6(sum_38_0_6, cout_38_0_6, sum_38_1_4, cout_37_0_5, sum_38_0_5);

wire sum_39_0_6, cout_39_0_6;

full_adder fa_39_0_6(sum_39_0_6, cout_39_0_6, sum_39_1_4, cout_38_0_5, sum_39_0_5);

wire sum_40_0_6, cout_40_0_6;

full_adder fa_40_0_6(sum_40_0_6, cout_40_0_6, sum_40_1_4, cout_39_0_5, sum_40_0_5);

wire sum_41_0_6, cout_41_0_6;

full_adder fa_41_0_6(sum_41_0_6, cout_41_0_6, sum_41_1_4, cout_40_0_5, sum_41_0_5);

wire sum_42_0_6, cout_42_0_6;

full_adder fa_42_0_6(sum_42_0_6, cout_42_0_6, sum_42_1_4, cout_41_0_5, sum_42_0_5);

wire sum_43_0_6, cout_43_0_6;

full_adder fa_43_0_6(sum_43_0_6, cout_43_0_6, sum_43_1_4, cout_42_0_5, sum_43_0_5);

wire sum_44_0_6, cout_44_0_6;

full_adder fa_44_0_6(sum_44_0_6, cout_44_0_6, sum_44_1_4, cout_43_0_5, sum_44_0_5);

wire sum_45_0_6, cout_45_0_6;

full_adder fa_45_0_6(sum_45_0_6, cout_45_0_6, sum_45_0_4, cout_44_0_5, sum_45_0_5);

wire sum_46_0_6, cout_46_0_6;

half_adder ha_46_0_6(sum_46_0_6, cout_46_0_6, cout_45_0_5, sum_46_0_5);

wire sum_47_0_6, cout_47_0_6;

half_adder ha_47_0_6(sum_47_0_6, cout_47_0_6, cout_46_0_5, sum_47_0_5);

wire sum_48_0_6, cout_48_0_6;

half_adder ha_48_0_6(sum_48_0_6, cout_48_0_6, cout_47_0_5, sum_48_0_5);

wire sum_49_0_6, cout_49_0_6;

half_adder ha_49_0_6(sum_49_0_6, cout_49_0_6, cout_48_0_5, sum_49_0_5);

wire sum_50_0_6, cout_50_0_6;

half_adder ha_50_0_6(sum_50_0_6, cout_50_0_6, cout_49_0_5, sum_50_0_5);

wire sum_51_0_6, cout_51_0_6;

half_adder ha_51_0_6(sum_51_0_6, cout_51_0_6, cout_50_0_5, sum_51_0_5);

wire sum_52_0_6, cout_52_0_6;

half_adder ha_52_0_6(sum_52_0_6, cout_52_0_6, cout_51_0_5, sum_52_0_5);

wire sum_53_0_6, cout_53_0_6;

half_adder ha_53_0_6(sum_53_0_6, cout_53_0_6, cout_52_0_5, sum_53_0_5);

wire sum_54_0_6, cout_54_0_6;

half_adder ha_54_0_6(sum_54_0_6, cout_54_0_6, cout_53_0_5, sum_54_0_5);

wire sum_55_0_6, cout_55_0_6;

half_adder ha_55_0_6(sum_55_0_6, cout_55_0_6, cout_54_0_5, sum_55_0_5);

wire sum_56_0_6, cout_56_0_6;

half_adder ha_56_0_6(sum_56_0_6, cout_56_0_6, cout_55_0_5, sum_56_0_5);

wire sum_57_0_6, cout_57_0_6;

half_adder ha_57_0_6(sum_57_0_6, cout_57_0_6, cout_56_0_5, sum_57_0_5);

wire sum_58_0_6, cout_58_0_6;

half_adder ha_58_0_6(sum_58_0_6, cout_58_0_6, cout_57_0_5, sum_58_0_5);

wire sum_59_0_6, cout_59_0_6;

half_adder ha_59_0_6(sum_59_0_6, cout_59_0_6, cout_58_0_5, sum_59_0_5);

wire sum_60_0_6, cout_60_0_6;

full_adder fa_60_0_6(sum_60_0_6, cout_60_0_6, cout_59_0_2, sum_60_0_2, cout_59_0_5);

wire sum_32_0_7, cout_32_0_7;

half_adder ha_32_0_7(sum_32_0_7, cout_32_0_7, sum_32_1_5, cout_31_0_6);

wire sum_33_0_7, cout_33_0_7;

full_adder fa_33_0_7(sum_33_0_7, cout_33_0_7, sum_33_1_5, cout_32_0_6, sum_33_0_6);

wire sum_34_0_7, cout_34_0_7;

full_adder fa_34_0_7(sum_34_0_7, cout_34_0_7, sum_34_1_5, cout_33_0_6, sum_34_0_6);

wire sum_35_0_7, cout_35_0_7;

full_adder fa_35_0_7(sum_35_0_7, cout_35_0_7, sum_35_1_5, cout_34_0_6, sum_35_0_6);

wire sum_36_0_7, cout_36_0_7;

full_adder fa_36_0_7(sum_36_0_7, cout_36_0_7, sum_36_1_5, cout_35_0_6, sum_36_0_6);

wire sum_37_0_7, cout_37_0_7;

full_adder fa_37_0_7(sum_37_0_7, cout_37_0_7, sum_37_0_5, cout_36_0_6, sum_37_0_6);

wire sum_38_0_7, cout_38_0_7;

half_adder ha_38_0_7(sum_38_0_7, cout_38_0_7, cout_37_0_6, sum_38_0_6);

wire sum_39_0_7, cout_39_0_7;

half_adder ha_39_0_7(sum_39_0_7, cout_39_0_7, cout_38_0_6, sum_39_0_6);

wire sum_40_0_7, cout_40_0_7;

half_adder ha_40_0_7(sum_40_0_7, cout_40_0_7, cout_39_0_6, sum_40_0_6);

wire sum_41_0_7, cout_41_0_7;

half_adder ha_41_0_7(sum_41_0_7, cout_41_0_7, cout_40_0_6, sum_41_0_6);

wire sum_42_0_7, cout_42_0_7;

half_adder ha_42_0_7(sum_42_0_7, cout_42_0_7, cout_41_0_6, sum_42_0_6);

wire sum_43_0_7, cout_43_0_7;

half_adder ha_43_0_7(sum_43_0_7, cout_43_0_7, cout_42_0_6, sum_43_0_6);

wire sum_44_0_7, cout_44_0_7;

half_adder ha_44_0_7(sum_44_0_7, cout_44_0_7, cout_43_0_6, sum_44_0_6);

wire sum_45_0_7, cout_45_0_7;

half_adder ha_45_0_7(sum_45_0_7, cout_45_0_7, cout_44_0_6, sum_45_0_6);

wire sum_46_0_7, cout_46_0_7;

half_adder ha_46_0_7(sum_46_0_7, cout_46_0_7, cout_45_0_6, sum_46_0_6);

wire sum_47_0_7, cout_47_0_7;

half_adder ha_47_0_7(sum_47_0_7, cout_47_0_7, cout_46_0_6, sum_47_0_6);

wire sum_48_0_7, cout_48_0_7;

half_adder ha_48_0_7(sum_48_0_7, cout_48_0_7, cout_47_0_6, sum_48_0_6);

wire sum_49_0_7, cout_49_0_7;

half_adder ha_49_0_7(sum_49_0_7, cout_49_0_7, cout_48_0_6, sum_49_0_6);

wire sum_50_0_7, cout_50_0_7;

half_adder ha_50_0_7(sum_50_0_7, cout_50_0_7, cout_49_0_6, sum_50_0_6);

wire sum_51_0_7, cout_51_0_7;

half_adder ha_51_0_7(sum_51_0_7, cout_51_0_7, cout_50_0_6, sum_51_0_6);

wire sum_52_0_7, cout_52_0_7;

half_adder ha_52_0_7(sum_52_0_7, cout_52_0_7, cout_51_0_6, sum_52_0_6);

wire sum_53_0_7, cout_53_0_7;

half_adder ha_53_0_7(sum_53_0_7, cout_53_0_7, cout_52_0_6, sum_53_0_6);

wire sum_54_0_7, cout_54_0_7;

half_adder ha_54_0_7(sum_54_0_7, cout_54_0_7, cout_53_0_6, sum_54_0_6);

wire sum_55_0_7, cout_55_0_7;

half_adder ha_55_0_7(sum_55_0_7, cout_55_0_7, cout_54_0_6, sum_55_0_6);

wire sum_56_0_7, cout_56_0_7;

half_adder ha_56_0_7(sum_56_0_7, cout_56_0_7, cout_55_0_6, sum_56_0_6);

wire sum_57_0_7, cout_57_0_7;

half_adder ha_57_0_7(sum_57_0_7, cout_57_0_7, cout_56_0_6, sum_57_0_6);

wire sum_58_0_7, cout_58_0_7;

half_adder ha_58_0_7(sum_58_0_7, cout_58_0_7, cout_57_0_6, sum_58_0_6);

wire sum_59_0_7, cout_59_0_7;

half_adder ha_59_0_7(sum_59_0_7, cout_59_0_7, cout_58_0_6, sum_59_0_6);

wire sum_60_0_7, cout_60_0_7;

half_adder ha_60_0_7(sum_60_0_7, cout_60_0_7, cout_59_0_6, sum_60_0_6);

wire sum_61_0_7, cout_61_0_7;

full_adder fa_61_0_7(sum_61_0_7, cout_61_0_7, cout_60_0_2, sum_61_0_2, cout_60_0_6);

wire sum_62_0_8, cout_62_0_8;

half_adder ha_62_0_8(sum_62_0_8, cout_62_0_8, A31B31, cout_61_0_2);

// ------------------------------------------------------------

// Adding using two CLA adders

wire [31:0] lsb_data_operandA, lsb_data_operandB;
wire lsb_cout;

assign lsb_data_operandA[31] = cout_30_0_6;
assign lsb_data_operandA[30] = cout_29_0_6;
assign lsb_data_operandA[29] = cout_28_0_6;
assign lsb_data_operandA[28] = cout_27_0_6;
assign lsb_data_operandA[27] = cout_26_0_6;
assign lsb_data_operandA[26] = cout_25_0_6;
assign lsb_data_operandA[25] = cout_24_0_6;
assign lsb_data_operandA[24] = cout_23_0_6;
assign lsb_data_operandA[23] = cout_22_0_6;
assign lsb_data_operandA[22] = sum_22_0_5;
assign lsb_data_operandA[21] = cout_20_0_5;
assign lsb_data_operandA[20] = cout_19_0_5;
assign lsb_data_operandA[19] = cout_18_0_5;
assign lsb_data_operandA[18] = cout_17_0_5;
assign lsb_data_operandA[17] = cout_16_0_5;
assign lsb_data_operandA[16] = cout_15_0_5;
assign lsb_data_operandA[15] = sum_15_0_4;
assign lsb_data_operandA[14] = cout_13_0_4;
assign lsb_data_operandA[13] = cout_12_0_4;
assign lsb_data_operandA[12] = cout_11_0_4;
assign lsb_data_operandA[11] = cout_10_0_4;
assign lsb_data_operandA[10] = sum_10_0_3;
assign lsb_data_operandA[9] = cout_8_0_3;
assign lsb_data_operandA[8] = cout_7_0_3;
assign lsb_data_operandA[7] = sum_7_0_2;
assign lsb_data_operandA[6] = cout_5_0_2;
assign lsb_data_operandA[5] = sum_5_0_1;
assign lsb_data_operandA[4] = cout_3_0_1;
assign lsb_data_operandA[3] = sum_3_0_0;
assign lsb_data_operandA[2] = A0B2;
assign lsb_data_operandA[1] = A1B0;
assign lsb_data_operandA[0] = A0B0;
// ------------------------------------------------------------

assign lsb_data_operandB[31] = sum_31_0_6;
assign lsb_data_operandB[30] = sum_30_0_6;
assign lsb_data_operandB[29] = sum_29_0_6;
assign lsb_data_operandB[28] = sum_28_0_6;
assign lsb_data_operandB[27] = sum_27_0_6;
assign lsb_data_operandB[26] = sum_26_0_6;
assign lsb_data_operandB[25] = sum_25_0_6;
assign lsb_data_operandB[24] = sum_24_0_6;
assign lsb_data_operandB[23] = sum_23_0_6;
assign lsb_data_operandB[22] = sum_22_0_6;
assign lsb_data_operandB[21] = sum_21_0_5;
assign lsb_data_operandB[20] = sum_20_0_5;
assign lsb_data_operandB[19] = sum_19_0_5;
assign lsb_data_operandB[18] = sum_18_0_5;
assign lsb_data_operandB[17] = sum_17_0_5;
assign lsb_data_operandB[16] = sum_16_0_5;
assign lsb_data_operandB[15] = sum_15_0_5;
assign lsb_data_operandB[14] = sum_14_0_4;
assign lsb_data_operandB[13] = sum_13_0_4;
assign lsb_data_operandB[12] = sum_12_0_4;
assign lsb_data_operandB[11] = sum_11_0_4;
assign lsb_data_operandB[10] = sum_10_0_4;
assign lsb_data_operandB[9] = sum_9_0_3;
assign lsb_data_operandB[8] = sum_8_0_3;
assign lsb_data_operandB[7] = sum_7_0_3;
assign lsb_data_operandB[6] = sum_6_0_2;
assign lsb_data_operandB[5] = sum_5_0_2;
assign lsb_data_operandB[4] = sum_4_0_1;
assign lsb_data_operandB[3] = sum_3_0_1;
assign lsb_data_operandB[2] = sum_2_0_0;
assign lsb_data_operandB[1] = A0B1;
assign lsb_data_operandB[0] = 1'b0;
cla_32 lsb_cla(data_result, lsb_cout, lsb_data_operandA, lsb_data_operandB, 1'b0);

// ------------------------------------------------------------

wire [31:0] msb_data_operandA, msb_data_operandB;
wire msb_cout;

assign msb_data_operandA[31] = cout_62_0_8;
assign msb_data_operandA[30] = cout_61_0_7;
assign msb_data_operandA[29] = cout_60_0_7;
assign msb_data_operandA[28] = cout_59_0_7;
assign msb_data_operandA[27] = cout_58_0_7;
assign msb_data_operandA[26] = cout_57_0_7;
assign msb_data_operandA[25] = cout_56_0_7;
assign msb_data_operandA[24] = cout_55_0_7;
assign msb_data_operandA[23] = cout_54_0_7;
assign msb_data_operandA[22] = cout_53_0_7;
assign msb_data_operandA[21] = cout_52_0_7;
assign msb_data_operandA[20] = cout_51_0_7;
assign msb_data_operandA[19] = cout_50_0_7;
assign msb_data_operandA[18] = cout_49_0_7;
assign msb_data_operandA[17] = cout_48_0_7;
assign msb_data_operandA[16] = cout_47_0_7;
assign msb_data_operandA[15] = cout_46_0_7;
assign msb_data_operandA[14] = cout_45_0_7;
assign msb_data_operandA[13] = cout_44_0_7;
assign msb_data_operandA[12] = cout_43_0_7;
assign msb_data_operandA[11] = cout_42_0_7;
assign msb_data_operandA[10] = cout_41_0_7;
assign msb_data_operandA[9] = cout_40_0_7;
assign msb_data_operandA[8] = cout_39_0_7;
assign msb_data_operandA[7] = cout_38_0_7;
assign msb_data_operandA[6] = cout_37_0_7;
assign msb_data_operandA[5] = cout_36_0_7;
assign msb_data_operandA[4] = cout_35_0_7;
assign msb_data_operandA[3] = cout_34_0_7;
assign msb_data_operandA[2] = cout_33_0_7;
assign msb_data_operandA[1] = cout_32_0_7;
assign msb_data_operandA[0] = sum_32_0_6;
// ------------------------------------------------------------

assign msb_data_operandB[31] = 1'b0;
assign msb_data_operandB[30] = sum_62_0_8;
assign msb_data_operandB[29] = sum_61_0_7;
assign msb_data_operandB[28] = sum_60_0_7;
assign msb_data_operandB[27] = sum_59_0_7;
assign msb_data_operandB[26] = sum_58_0_7;
assign msb_data_operandB[25] = sum_57_0_7;
assign msb_data_operandB[24] = sum_56_0_7;
assign msb_data_operandB[23] = sum_55_0_7;
assign msb_data_operandB[22] = sum_54_0_7;
assign msb_data_operandB[21] = sum_53_0_7;
assign msb_data_operandB[20] = sum_52_0_7;
assign msb_data_operandB[19] = sum_51_0_7;
assign msb_data_operandB[18] = sum_50_0_7;
assign msb_data_operandB[17] = sum_49_0_7;
assign msb_data_operandB[16] = sum_48_0_7;
assign msb_data_operandB[15] = sum_47_0_7;
assign msb_data_operandB[14] = sum_46_0_7;
assign msb_data_operandB[13] = sum_45_0_7;
assign msb_data_operandB[12] = sum_44_0_7;
assign msb_data_operandB[11] = sum_43_0_7;
assign msb_data_operandB[10] = sum_42_0_7;
assign msb_data_operandB[9] = sum_41_0_7;
assign msb_data_operandB[8] = sum_40_0_7;
assign msb_data_operandB[7] = sum_39_0_7;
assign msb_data_operandB[6] = sum_38_0_7;
assign msb_data_operandB[5] = sum_37_0_7;
assign msb_data_operandB[4] = sum_36_0_7;
assign msb_data_operandB[3] = sum_35_0_7;
assign msb_data_operandB[2] = sum_34_0_7;
assign msb_data_operandB[1] = sum_33_0_7;
assign msb_data_operandB[0] = sum_32_0_7;
cla_32 msb_cla(msb_data_result, msb_cout, msb_data_operandA, msb_data_operandB, lsb_cout);

// ------------------------------------------------------------

// Check for overflow by checking whether all msb 33 bits are the same
wire and_result, nor_result;
and and_overflow(and_result, msb_data_result[31], msb_data_result[30], msb_data_result[29], msb_data_result[28], msb_data_result[27], msb_data_result[26], msb_data_result[25], msb_data_result[24], msb_data_result[23], msb_data_result[22], msb_data_result[21], msb_data_result[20], msb_data_result[19], msb_data_result[18], msb_data_result[17], msb_data_result[16], msb_data_result[15], msb_data_result[14], msb_data_result[13], msb_data_result[12], msb_data_result[11], msb_data_result[10], msb_data_result[9], msb_data_result[8], msb_data_result[7], msb_data_result[6], msb_data_result[5], msb_data_result[4], msb_data_result[3], msb_data_result[2], msb_data_result[1], msb_data_result[0], data_result[31]);

nor nor_overflow(nor_result, msb_data_result[31], msb_data_result[30], msb_data_result[29], msb_data_result[28], msb_data_result[27], msb_data_result[26], msb_data_result[25], msb_data_result[24], msb_data_result[23], msb_data_result[22], msb_data_result[21], msb_data_result[20], msb_data_result[19], msb_data_result[18], msb_data_result[17], msb_data_result[16], msb_data_result[15], msb_data_result[14], msb_data_result[13], msb_data_result[12], msb_data_result[11], msb_data_result[10], msb_data_result[9], msb_data_result[8], msb_data_result[7], msb_data_result[6], msb_data_result[5], msb_data_result[4], msb_data_result[3], msb_data_result[2], msb_data_result[1], msb_data_result[0], data_result[31]);

xnor exception(data_exception, and_result, nor_result);
endmodule
module multdiv(
	data_operandA, data_operandB, 
	ctrl_MULT, ctrl_DIV, 
	clock, 
	data_result, data_exception, data_resultRDY);

    input [31:0] data_operandA, data_operandB;
    input ctrl_MULT, ctrl_DIV, clock;

    output [31:0] data_result;
    output data_exception, data_resultRDY;

    // add your code here
    wire [31:0] mult_result, div_result;
    multiplier mult(mult_result, data_resultRDY, data_exception, data_operandA, data_operandB, clock);
    // divider div(div_result, data_resultRDY, data_exception, data_operandA, data_operandB, clock);

    assign data_result = mult_result;
endmodule